/home/linux/ieng6/ee260bwi25/ttalapaneni/ECE260B_course_project/Git_organized_folder/ECE260B_course_project/pnr/part3_hier/pnr_2_SRAM_V3/subckt/sram_w16.lef