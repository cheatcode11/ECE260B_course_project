##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Tue Mar  4 02:09:13 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 461.8000 BY 459.2000 ;
  FOREIGN fullchip 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 54.9500 0.6000 55.0500 ;
    END
  END clk
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 218.9500 0.6000 219.0500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 216.9500 0.6000 217.0500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 214.9500 0.6000 215.0500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 212.9500 0.6000 213.0500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 210.9500 0.6000 211.0500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 208.9500 0.6000 209.0500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 206.9500 0.6000 207.0500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 204.9500 0.6000 205.0500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 202.9500 0.6000 203.0500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 200.9500 0.6000 201.0500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 198.9500 0.6000 199.0500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 196.9500 0.6000 197.0500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 194.9500 0.6000 195.0500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 192.9500 0.6000 193.0500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 190.9500 0.6000 191.0500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 188.9500 0.6000 189.0500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 186.9500 0.6000 187.0500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 184.9500 0.6000 185.0500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 182.9500 0.6000 183.0500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 180.9500 0.6000 181.0500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 178.9500 0.6000 179.0500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 176.9500 0.6000 177.0500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 174.9500 0.6000 175.0500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 172.9500 0.6000 173.0500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 170.9500 0.6000 171.0500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 168.9500 0.6000 169.0500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 166.9500 0.6000 167.0500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 164.9500 0.6000 165.0500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 162.9500 0.6000 163.0500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 160.9500 0.6000 161.0500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 158.9500 0.6000 159.0500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 156.9500 0.6000 157.0500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 154.9500 0.6000 155.0500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 152.9500 0.6000 153.0500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 150.9500 0.6000 151.0500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 148.9500 0.6000 149.0500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 146.9500 0.6000 147.0500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 144.9500 0.6000 145.0500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 142.9500 0.6000 143.0500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 140.9500 0.6000 141.0500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 138.9500 0.6000 139.0500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 136.9500 0.6000 137.0500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 134.9500 0.6000 135.0500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 132.9500 0.6000 133.0500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 130.9500 0.6000 131.0500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 128.9500 0.6000 129.0500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 126.9500 0.6000 127.0500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 124.9500 0.6000 125.0500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 122.9500 0.6000 123.0500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 120.9500 0.6000 121.0500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 118.9500 0.6000 119.0500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 116.9500 0.6000 117.0500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 114.9500 0.6000 115.0500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 112.9500 0.6000 113.0500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 110.9500 0.6000 111.0500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 108.9500 0.6000 109.0500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 106.9500 0.6000 107.0500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 104.9500 0.6000 105.0500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 102.9500 0.6000 103.0500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 100.9500 0.6000 101.0500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 98.9500 0.6000 99.0500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 96.9500 0.6000 97.0500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 94.9500 0.6000 95.0500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 92.9500 0.6000 93.0500 ;
    END
  END mem_in[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 88.9500 0.6000 89.0500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 86.9500 0.6000 87.0500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 84.9500 0.6000 85.0500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 82.9500 0.6000 83.0500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 80.9500 0.6000 81.0500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 78.9500 0.6000 79.0500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 76.9500 0.6000 77.0500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 74.9500 0.6000 75.0500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 72.9500 0.6000 73.0500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 70.9500 0.6000 71.0500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 68.9500 0.6000 69.0500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 66.9500 0.6000 67.0500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 64.9500 0.6000 65.0500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 62.9500 0.6000 63.0500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 60.9500 0.6000 61.0500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 58.9500 0.6000 59.0500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 56.9500 0.6000 57.0500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 90.9500 0.6000 91.0500 ;
    END
  END reset
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 373.0500 0.0000 373.1500 0.6000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.0500 0.0000 371.1500 0.6000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.0500 0.0000 369.1500 0.6000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.0500 0.0000 367.1500 0.6000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 365.0500 0.0000 365.1500 0.6000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.0500 0.0000 363.1500 0.6000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.0500 0.0000 361.1500 0.6000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.0500 0.0000 359.1500 0.6000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.0500 0.0000 357.1500 0.6000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.0500 0.0000 355.1500 0.6000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.0500 0.0000 353.1500 0.6000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.0500 0.0000 351.1500 0.6000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.0500 0.0000 349.1500 0.6000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.0500 0.0000 347.1500 0.6000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.0500 0.0000 345.1500 0.6000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.0500 0.0000 343.1500 0.6000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.0500 0.0000 341.1500 0.6000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.0500 0.0000 339.1500 0.6000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.0500 0.0000 337.1500 0.6000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.0500 0.0000 335.1500 0.6000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.0500 0.0000 333.1500 0.6000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.0500 0.0000 331.1500 0.6000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.0500 0.0000 329.1500 0.6000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.0500 0.0000 327.1500 0.6000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.0500 0.0000 325.1500 0.6000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.0500 0.0000 323.1500 0.6000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.0500 0.0000 321.1500 0.6000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.0500 0.0000 319.1500 0.6000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.0500 0.0000 317.1500 0.6000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.0500 0.0000 315.1500 0.6000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.0500 0.0000 313.1500 0.6000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.0500 0.0000 311.1500 0.6000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.0500 0.0000 309.1500 0.6000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.0500 0.0000 307.1500 0.6000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 305.0500 0.0000 305.1500 0.6000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.0500 0.0000 303.1500 0.6000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 301.0500 0.0000 301.1500 0.6000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 299.0500 0.0000 299.1500 0.6000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 297.0500 0.0000 297.1500 0.6000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.0500 0.0000 295.1500 0.6000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 293.0500 0.0000 293.1500 0.6000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.0500 0.0000 291.1500 0.6000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 289.0500 0.0000 289.1500 0.6000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 287.0500 0.0000 287.1500 0.6000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 285.0500 0.0000 285.1500 0.6000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 283.0500 0.0000 283.1500 0.6000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 281.0500 0.0000 281.1500 0.6000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 279.0500 0.0000 279.1500 0.6000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.0500 0.0000 277.1500 0.6000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 275.0500 0.0000 275.1500 0.6000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.0500 0.0000 273.1500 0.6000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 271.0500 0.0000 271.1500 0.6000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 269.0500 0.0000 269.1500 0.6000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.0500 0.0000 267.1500 0.6000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 265.0500 0.0000 265.1500 0.6000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 263.0500 0.0000 263.1500 0.6000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 261.0500 0.0000 261.1500 0.6000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.0500 0.0000 259.1500 0.6000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 257.0500 0.0000 257.1500 0.6000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.0500 0.0000 255.1500 0.6000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 253.0500 0.0000 253.1500 0.6000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 251.0500 0.0000 251.1500 0.6000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 249.0500 0.0000 249.1500 0.6000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.0500 0.0000 247.1500 0.6000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 245.0500 0.0000 245.1500 0.6000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.0500 0.0000 243.1500 0.6000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.0500 0.0000 241.1500 0.6000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 239.0500 0.0000 239.1500 0.6000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.0500 0.0000 237.1500 0.6000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.0500 0.0000 235.1500 0.6000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.0500 0.0000 233.1500 0.6000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.0500 0.0000 231.1500 0.6000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 229.0500 0.0000 229.1500 0.6000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.0500 0.0000 227.1500 0.6000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 225.0500 0.0000 225.1500 0.6000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.0500 0.0000 223.1500 0.6000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 221.0500 0.0000 221.1500 0.6000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.0500 0.0000 219.1500 0.6000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.0500 0.0000 217.1500 0.6000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.0500 0.0000 215.1500 0.6000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.0500 0.0000 213.1500 0.6000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.0500 0.0000 211.1500 0.6000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.0500 0.0000 209.1500 0.6000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.0500 0.0000 207.1500 0.6000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.0500 0.0000 205.1500 0.6000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.0500 0.0000 203.1500 0.6000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.0500 0.0000 201.1500 0.6000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.0500 0.0000 199.1500 0.6000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.0500 0.0000 197.1500 0.6000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.0500 0.0000 195.1500 0.6000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.0500 0.0000 193.1500 0.6000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.0500 0.0000 191.1500 0.6000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.0500 0.0000 189.1500 0.6000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.0500 0.0000 187.1500 0.6000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 185.0500 0.0000 185.1500 0.6000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.0500 0.0000 183.1500 0.6000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.0500 0.0000 181.1500 0.6000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.0500 0.0000 179.1500 0.6000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.0500 0.0000 177.1500 0.6000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.0500 0.0000 175.1500 0.6000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.0500 0.0000 173.1500 0.6000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.0500 0.0000 171.1500 0.6000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.0500 0.0000 169.1500 0.6000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.0500 0.0000 167.1500 0.6000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.0500 0.0000 165.1500 0.6000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.0500 0.0000 163.1500 0.6000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.0500 0.0000 161.1500 0.6000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.0500 0.0000 159.1500 0.6000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.0500 0.0000 157.1500 0.6000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.0500 0.0000 155.1500 0.6000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.0500 0.0000 153.1500 0.6000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.0500 0.0000 151.1500 0.6000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.0500 0.0000 149.1500 0.6000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.0500 0.0000 147.1500 0.6000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.0500 0.0000 145.1500 0.6000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.0500 0.0000 143.1500 0.6000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.0500 0.0000 141.1500 0.6000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.0500 0.0000 139.1500 0.6000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.0500 0.0000 137.1500 0.6000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.0500 0.0000 135.1500 0.6000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.0500 0.0000 133.1500 0.6000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.0500 0.0000 131.1500 0.6000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.0500 0.0000 129.1500 0.6000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.0500 0.0000 127.1500 0.6000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.0500 0.0000 125.1500 0.6000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.0500 0.0000 123.1500 0.6000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.0500 0.0000 121.1500 0.6000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.0500 0.0000 119.1500 0.6000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.0500 0.0000 117.1500 0.6000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.0500 0.0000 115.1500 0.6000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.0500 0.0000 113.1500 0.6000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.0500 0.0000 111.1500 0.6000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.0500 0.0000 109.1500 0.6000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.0500 0.0000 107.1500 0.6000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.0500 0.0000 105.1500 0.6000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.0500 0.0000 103.1500 0.6000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.0500 0.0000 101.1500 0.6000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.0500 0.0000 99.1500 0.6000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.0500 0.0000 97.1500 0.6000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.0500 0.0000 95.1500 0.6000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.0500 0.0000 93.1500 0.6000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.0500 0.0000 91.1500 0.6000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.0500 0.0000 89.1500 0.6000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.0500 0.0000 87.1500 0.6000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.0500 0.0000 85.1500 0.6000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.0500 0.0000 83.1500 0.6000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.0500 0.0000 81.1500 0.6000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.0500 0.0000 79.1500 0.6000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.0500 0.0000 77.1500 0.6000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.0500 0.0000 75.1500 0.6000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.0500 0.0000 73.1500 0.6000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.0500 0.0000 71.1500 0.6000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.0500 0.0000 69.1500 0.6000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.0500 0.0000 67.1500 0.6000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.0500 0.0000 65.1500 0.6000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.0500 0.0000 63.1500 0.6000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.0500 0.0000 61.1500 0.6000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.0500 0.0000 59.1500 0.6000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.0500 0.0000 57.1500 0.6000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.0500 0.0000 55.1500 0.6000 ;
    END
  END out[0]
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 461.8000 459.2000 ;
    LAYER M2 ;
      RECT 0.0000 0.7000 461.8000 459.2000 ;
      RECT 373.2500 0.0000 461.8000 0.7000 ;
      RECT 371.2500 0.0000 372.9500 0.7000 ;
      RECT 369.2500 0.0000 370.9500 0.7000 ;
      RECT 367.2500 0.0000 368.9500 0.7000 ;
      RECT 365.2500 0.0000 366.9500 0.7000 ;
      RECT 363.2500 0.0000 364.9500 0.7000 ;
      RECT 361.2500 0.0000 362.9500 0.7000 ;
      RECT 359.2500 0.0000 360.9500 0.7000 ;
      RECT 357.2500 0.0000 358.9500 0.7000 ;
      RECT 355.2500 0.0000 356.9500 0.7000 ;
      RECT 353.2500 0.0000 354.9500 0.7000 ;
      RECT 351.2500 0.0000 352.9500 0.7000 ;
      RECT 349.2500 0.0000 350.9500 0.7000 ;
      RECT 347.2500 0.0000 348.9500 0.7000 ;
      RECT 345.2500 0.0000 346.9500 0.7000 ;
      RECT 343.2500 0.0000 344.9500 0.7000 ;
      RECT 341.2500 0.0000 342.9500 0.7000 ;
      RECT 339.2500 0.0000 340.9500 0.7000 ;
      RECT 337.2500 0.0000 338.9500 0.7000 ;
      RECT 335.2500 0.0000 336.9500 0.7000 ;
      RECT 333.2500 0.0000 334.9500 0.7000 ;
      RECT 331.2500 0.0000 332.9500 0.7000 ;
      RECT 329.2500 0.0000 330.9500 0.7000 ;
      RECT 327.2500 0.0000 328.9500 0.7000 ;
      RECT 325.2500 0.0000 326.9500 0.7000 ;
      RECT 323.2500 0.0000 324.9500 0.7000 ;
      RECT 321.2500 0.0000 322.9500 0.7000 ;
      RECT 319.2500 0.0000 320.9500 0.7000 ;
      RECT 317.2500 0.0000 318.9500 0.7000 ;
      RECT 315.2500 0.0000 316.9500 0.7000 ;
      RECT 313.2500 0.0000 314.9500 0.7000 ;
      RECT 311.2500 0.0000 312.9500 0.7000 ;
      RECT 309.2500 0.0000 310.9500 0.7000 ;
      RECT 307.2500 0.0000 308.9500 0.7000 ;
      RECT 305.2500 0.0000 306.9500 0.7000 ;
      RECT 303.2500 0.0000 304.9500 0.7000 ;
      RECT 301.2500 0.0000 302.9500 0.7000 ;
      RECT 299.2500 0.0000 300.9500 0.7000 ;
      RECT 297.2500 0.0000 298.9500 0.7000 ;
      RECT 295.2500 0.0000 296.9500 0.7000 ;
      RECT 293.2500 0.0000 294.9500 0.7000 ;
      RECT 291.2500 0.0000 292.9500 0.7000 ;
      RECT 289.2500 0.0000 290.9500 0.7000 ;
      RECT 287.2500 0.0000 288.9500 0.7000 ;
      RECT 285.2500 0.0000 286.9500 0.7000 ;
      RECT 283.2500 0.0000 284.9500 0.7000 ;
      RECT 281.2500 0.0000 282.9500 0.7000 ;
      RECT 279.2500 0.0000 280.9500 0.7000 ;
      RECT 277.2500 0.0000 278.9500 0.7000 ;
      RECT 275.2500 0.0000 276.9500 0.7000 ;
      RECT 273.2500 0.0000 274.9500 0.7000 ;
      RECT 271.2500 0.0000 272.9500 0.7000 ;
      RECT 269.2500 0.0000 270.9500 0.7000 ;
      RECT 267.2500 0.0000 268.9500 0.7000 ;
      RECT 265.2500 0.0000 266.9500 0.7000 ;
      RECT 263.2500 0.0000 264.9500 0.7000 ;
      RECT 261.2500 0.0000 262.9500 0.7000 ;
      RECT 259.2500 0.0000 260.9500 0.7000 ;
      RECT 257.2500 0.0000 258.9500 0.7000 ;
      RECT 255.2500 0.0000 256.9500 0.7000 ;
      RECT 253.2500 0.0000 254.9500 0.7000 ;
      RECT 251.2500 0.0000 252.9500 0.7000 ;
      RECT 249.2500 0.0000 250.9500 0.7000 ;
      RECT 247.2500 0.0000 248.9500 0.7000 ;
      RECT 245.2500 0.0000 246.9500 0.7000 ;
      RECT 243.2500 0.0000 244.9500 0.7000 ;
      RECT 241.2500 0.0000 242.9500 0.7000 ;
      RECT 239.2500 0.0000 240.9500 0.7000 ;
      RECT 237.2500 0.0000 238.9500 0.7000 ;
      RECT 235.2500 0.0000 236.9500 0.7000 ;
      RECT 233.2500 0.0000 234.9500 0.7000 ;
      RECT 231.2500 0.0000 232.9500 0.7000 ;
      RECT 229.2500 0.0000 230.9500 0.7000 ;
      RECT 227.2500 0.0000 228.9500 0.7000 ;
      RECT 225.2500 0.0000 226.9500 0.7000 ;
      RECT 223.2500 0.0000 224.9500 0.7000 ;
      RECT 221.2500 0.0000 222.9500 0.7000 ;
      RECT 219.2500 0.0000 220.9500 0.7000 ;
      RECT 217.2500 0.0000 218.9500 0.7000 ;
      RECT 215.2500 0.0000 216.9500 0.7000 ;
      RECT 213.2500 0.0000 214.9500 0.7000 ;
      RECT 211.2500 0.0000 212.9500 0.7000 ;
      RECT 209.2500 0.0000 210.9500 0.7000 ;
      RECT 207.2500 0.0000 208.9500 0.7000 ;
      RECT 205.2500 0.0000 206.9500 0.7000 ;
      RECT 203.2500 0.0000 204.9500 0.7000 ;
      RECT 201.2500 0.0000 202.9500 0.7000 ;
      RECT 199.2500 0.0000 200.9500 0.7000 ;
      RECT 197.2500 0.0000 198.9500 0.7000 ;
      RECT 195.2500 0.0000 196.9500 0.7000 ;
      RECT 193.2500 0.0000 194.9500 0.7000 ;
      RECT 191.2500 0.0000 192.9500 0.7000 ;
      RECT 189.2500 0.0000 190.9500 0.7000 ;
      RECT 187.2500 0.0000 188.9500 0.7000 ;
      RECT 185.2500 0.0000 186.9500 0.7000 ;
      RECT 183.2500 0.0000 184.9500 0.7000 ;
      RECT 181.2500 0.0000 182.9500 0.7000 ;
      RECT 179.2500 0.0000 180.9500 0.7000 ;
      RECT 177.2500 0.0000 178.9500 0.7000 ;
      RECT 175.2500 0.0000 176.9500 0.7000 ;
      RECT 173.2500 0.0000 174.9500 0.7000 ;
      RECT 171.2500 0.0000 172.9500 0.7000 ;
      RECT 169.2500 0.0000 170.9500 0.7000 ;
      RECT 167.2500 0.0000 168.9500 0.7000 ;
      RECT 165.2500 0.0000 166.9500 0.7000 ;
      RECT 163.2500 0.0000 164.9500 0.7000 ;
      RECT 161.2500 0.0000 162.9500 0.7000 ;
      RECT 159.2500 0.0000 160.9500 0.7000 ;
      RECT 157.2500 0.0000 158.9500 0.7000 ;
      RECT 155.2500 0.0000 156.9500 0.7000 ;
      RECT 153.2500 0.0000 154.9500 0.7000 ;
      RECT 151.2500 0.0000 152.9500 0.7000 ;
      RECT 149.2500 0.0000 150.9500 0.7000 ;
      RECT 147.2500 0.0000 148.9500 0.7000 ;
      RECT 145.2500 0.0000 146.9500 0.7000 ;
      RECT 143.2500 0.0000 144.9500 0.7000 ;
      RECT 141.2500 0.0000 142.9500 0.7000 ;
      RECT 139.2500 0.0000 140.9500 0.7000 ;
      RECT 137.2500 0.0000 138.9500 0.7000 ;
      RECT 135.2500 0.0000 136.9500 0.7000 ;
      RECT 133.2500 0.0000 134.9500 0.7000 ;
      RECT 131.2500 0.0000 132.9500 0.7000 ;
      RECT 129.2500 0.0000 130.9500 0.7000 ;
      RECT 127.2500 0.0000 128.9500 0.7000 ;
      RECT 125.2500 0.0000 126.9500 0.7000 ;
      RECT 123.2500 0.0000 124.9500 0.7000 ;
      RECT 121.2500 0.0000 122.9500 0.7000 ;
      RECT 119.2500 0.0000 120.9500 0.7000 ;
      RECT 117.2500 0.0000 118.9500 0.7000 ;
      RECT 115.2500 0.0000 116.9500 0.7000 ;
      RECT 113.2500 0.0000 114.9500 0.7000 ;
      RECT 111.2500 0.0000 112.9500 0.7000 ;
      RECT 109.2500 0.0000 110.9500 0.7000 ;
      RECT 107.2500 0.0000 108.9500 0.7000 ;
      RECT 105.2500 0.0000 106.9500 0.7000 ;
      RECT 103.2500 0.0000 104.9500 0.7000 ;
      RECT 101.2500 0.0000 102.9500 0.7000 ;
      RECT 99.2500 0.0000 100.9500 0.7000 ;
      RECT 97.2500 0.0000 98.9500 0.7000 ;
      RECT 95.2500 0.0000 96.9500 0.7000 ;
      RECT 93.2500 0.0000 94.9500 0.7000 ;
      RECT 91.2500 0.0000 92.9500 0.7000 ;
      RECT 89.2500 0.0000 90.9500 0.7000 ;
      RECT 87.2500 0.0000 88.9500 0.7000 ;
      RECT 85.2500 0.0000 86.9500 0.7000 ;
      RECT 83.2500 0.0000 84.9500 0.7000 ;
      RECT 81.2500 0.0000 82.9500 0.7000 ;
      RECT 79.2500 0.0000 80.9500 0.7000 ;
      RECT 77.2500 0.0000 78.9500 0.7000 ;
      RECT 75.2500 0.0000 76.9500 0.7000 ;
      RECT 73.2500 0.0000 74.9500 0.7000 ;
      RECT 71.2500 0.0000 72.9500 0.7000 ;
      RECT 69.2500 0.0000 70.9500 0.7000 ;
      RECT 67.2500 0.0000 68.9500 0.7000 ;
      RECT 65.2500 0.0000 66.9500 0.7000 ;
      RECT 63.2500 0.0000 64.9500 0.7000 ;
      RECT 61.2500 0.0000 62.9500 0.7000 ;
      RECT 59.2500 0.0000 60.9500 0.7000 ;
      RECT 57.2500 0.0000 58.9500 0.7000 ;
      RECT 55.2500 0.0000 56.9500 0.7000 ;
      RECT 0.0000 0.0000 54.9500 0.7000 ;
    LAYER M3 ;
      RECT 0.0000 219.1500 461.8000 459.2000 ;
      RECT 0.7000 218.8500 461.8000 219.1500 ;
      RECT 0.0000 217.1500 461.8000 218.8500 ;
      RECT 0.7000 216.8500 461.8000 217.1500 ;
      RECT 0.0000 215.1500 461.8000 216.8500 ;
      RECT 0.7000 214.8500 461.8000 215.1500 ;
      RECT 0.0000 213.1500 461.8000 214.8500 ;
      RECT 0.7000 212.8500 461.8000 213.1500 ;
      RECT 0.0000 211.1500 461.8000 212.8500 ;
      RECT 0.7000 210.8500 461.8000 211.1500 ;
      RECT 0.0000 209.1500 461.8000 210.8500 ;
      RECT 0.7000 208.8500 461.8000 209.1500 ;
      RECT 0.0000 207.1500 461.8000 208.8500 ;
      RECT 0.7000 206.8500 461.8000 207.1500 ;
      RECT 0.0000 205.1500 461.8000 206.8500 ;
      RECT 0.7000 204.8500 461.8000 205.1500 ;
      RECT 0.0000 203.1500 461.8000 204.8500 ;
      RECT 0.7000 202.8500 461.8000 203.1500 ;
      RECT 0.0000 201.1500 461.8000 202.8500 ;
      RECT 0.7000 200.8500 461.8000 201.1500 ;
      RECT 0.0000 199.1500 461.8000 200.8500 ;
      RECT 0.7000 198.8500 461.8000 199.1500 ;
      RECT 0.0000 197.1500 461.8000 198.8500 ;
      RECT 0.7000 196.8500 461.8000 197.1500 ;
      RECT 0.0000 195.1500 461.8000 196.8500 ;
      RECT 0.7000 194.8500 461.8000 195.1500 ;
      RECT 0.0000 193.1500 461.8000 194.8500 ;
      RECT 0.7000 192.8500 461.8000 193.1500 ;
      RECT 0.0000 191.1500 461.8000 192.8500 ;
      RECT 0.7000 190.8500 461.8000 191.1500 ;
      RECT 0.0000 189.1500 461.8000 190.8500 ;
      RECT 0.7000 188.8500 461.8000 189.1500 ;
      RECT 0.0000 187.1500 461.8000 188.8500 ;
      RECT 0.7000 186.8500 461.8000 187.1500 ;
      RECT 0.0000 185.1500 461.8000 186.8500 ;
      RECT 0.7000 184.8500 461.8000 185.1500 ;
      RECT 0.0000 183.1500 461.8000 184.8500 ;
      RECT 0.7000 182.8500 461.8000 183.1500 ;
      RECT 0.0000 181.1500 461.8000 182.8500 ;
      RECT 0.7000 180.8500 461.8000 181.1500 ;
      RECT 0.0000 179.1500 461.8000 180.8500 ;
      RECT 0.7000 178.8500 461.8000 179.1500 ;
      RECT 0.0000 177.1500 461.8000 178.8500 ;
      RECT 0.7000 176.8500 461.8000 177.1500 ;
      RECT 0.0000 175.1500 461.8000 176.8500 ;
      RECT 0.7000 174.8500 461.8000 175.1500 ;
      RECT 0.0000 173.1500 461.8000 174.8500 ;
      RECT 0.7000 172.8500 461.8000 173.1500 ;
      RECT 0.0000 171.1500 461.8000 172.8500 ;
      RECT 0.7000 170.8500 461.8000 171.1500 ;
      RECT 0.0000 169.1500 461.8000 170.8500 ;
      RECT 0.7000 168.8500 461.8000 169.1500 ;
      RECT 0.0000 167.1500 461.8000 168.8500 ;
      RECT 0.7000 166.8500 461.8000 167.1500 ;
      RECT 0.0000 165.1500 461.8000 166.8500 ;
      RECT 0.7000 164.8500 461.8000 165.1500 ;
      RECT 0.0000 163.1500 461.8000 164.8500 ;
      RECT 0.7000 162.8500 461.8000 163.1500 ;
      RECT 0.0000 161.1500 461.8000 162.8500 ;
      RECT 0.7000 160.8500 461.8000 161.1500 ;
      RECT 0.0000 159.1500 461.8000 160.8500 ;
      RECT 0.7000 158.8500 461.8000 159.1500 ;
      RECT 0.0000 157.1500 461.8000 158.8500 ;
      RECT 0.7000 156.8500 461.8000 157.1500 ;
      RECT 0.0000 155.1500 461.8000 156.8500 ;
      RECT 0.7000 154.8500 461.8000 155.1500 ;
      RECT 0.0000 153.1500 461.8000 154.8500 ;
      RECT 0.7000 152.8500 461.8000 153.1500 ;
      RECT 0.0000 151.1500 461.8000 152.8500 ;
      RECT 0.7000 150.8500 461.8000 151.1500 ;
      RECT 0.0000 149.1500 461.8000 150.8500 ;
      RECT 0.7000 148.8500 461.8000 149.1500 ;
      RECT 0.0000 147.1500 461.8000 148.8500 ;
      RECT 0.7000 146.8500 461.8000 147.1500 ;
      RECT 0.0000 145.1500 461.8000 146.8500 ;
      RECT 0.7000 144.8500 461.8000 145.1500 ;
      RECT 0.0000 143.1500 461.8000 144.8500 ;
      RECT 0.7000 142.8500 461.8000 143.1500 ;
      RECT 0.0000 141.1500 461.8000 142.8500 ;
      RECT 0.7000 140.8500 461.8000 141.1500 ;
      RECT 0.0000 139.1500 461.8000 140.8500 ;
      RECT 0.7000 138.8500 461.8000 139.1500 ;
      RECT 0.0000 137.1500 461.8000 138.8500 ;
      RECT 0.7000 136.8500 461.8000 137.1500 ;
      RECT 0.0000 135.1500 461.8000 136.8500 ;
      RECT 0.7000 134.8500 461.8000 135.1500 ;
      RECT 0.0000 133.1500 461.8000 134.8500 ;
      RECT 0.7000 132.8500 461.8000 133.1500 ;
      RECT 0.0000 131.1500 461.8000 132.8500 ;
      RECT 0.7000 130.8500 461.8000 131.1500 ;
      RECT 0.0000 129.1500 461.8000 130.8500 ;
      RECT 0.7000 128.8500 461.8000 129.1500 ;
      RECT 0.0000 127.1500 461.8000 128.8500 ;
      RECT 0.7000 126.8500 461.8000 127.1500 ;
      RECT 0.0000 125.1500 461.8000 126.8500 ;
      RECT 0.7000 124.8500 461.8000 125.1500 ;
      RECT 0.0000 123.1500 461.8000 124.8500 ;
      RECT 0.7000 122.8500 461.8000 123.1500 ;
      RECT 0.0000 121.1500 461.8000 122.8500 ;
      RECT 0.7000 120.8500 461.8000 121.1500 ;
      RECT 0.0000 119.1500 461.8000 120.8500 ;
      RECT 0.7000 118.8500 461.8000 119.1500 ;
      RECT 0.0000 117.1500 461.8000 118.8500 ;
      RECT 0.7000 116.8500 461.8000 117.1500 ;
      RECT 0.0000 115.1500 461.8000 116.8500 ;
      RECT 0.7000 114.8500 461.8000 115.1500 ;
      RECT 0.0000 113.1500 461.8000 114.8500 ;
      RECT 0.7000 112.8500 461.8000 113.1500 ;
      RECT 0.0000 111.1500 461.8000 112.8500 ;
      RECT 0.7000 110.8500 461.8000 111.1500 ;
      RECT 0.0000 109.1500 461.8000 110.8500 ;
      RECT 0.7000 108.8500 461.8000 109.1500 ;
      RECT 0.0000 107.1500 461.8000 108.8500 ;
      RECT 0.7000 106.8500 461.8000 107.1500 ;
      RECT 0.0000 105.1500 461.8000 106.8500 ;
      RECT 0.7000 104.8500 461.8000 105.1500 ;
      RECT 0.0000 103.1500 461.8000 104.8500 ;
      RECT 0.7000 102.8500 461.8000 103.1500 ;
      RECT 0.0000 101.1500 461.8000 102.8500 ;
      RECT 0.7000 100.8500 461.8000 101.1500 ;
      RECT 0.0000 99.1500 461.8000 100.8500 ;
      RECT 0.7000 98.8500 461.8000 99.1500 ;
      RECT 0.0000 97.1500 461.8000 98.8500 ;
      RECT 0.7000 96.8500 461.8000 97.1500 ;
      RECT 0.0000 95.1500 461.8000 96.8500 ;
      RECT 0.7000 94.8500 461.8000 95.1500 ;
      RECT 0.0000 93.1500 461.8000 94.8500 ;
      RECT 0.7000 92.8500 461.8000 93.1500 ;
      RECT 0.0000 91.1500 461.8000 92.8500 ;
      RECT 0.7000 90.8500 461.8000 91.1500 ;
      RECT 0.0000 89.1500 461.8000 90.8500 ;
      RECT 0.7000 88.8500 461.8000 89.1500 ;
      RECT 0.0000 87.1500 461.8000 88.8500 ;
      RECT 0.7000 86.8500 461.8000 87.1500 ;
      RECT 0.0000 85.1500 461.8000 86.8500 ;
      RECT 0.7000 84.8500 461.8000 85.1500 ;
      RECT 0.0000 83.1500 461.8000 84.8500 ;
      RECT 0.7000 82.8500 461.8000 83.1500 ;
      RECT 0.0000 81.1500 461.8000 82.8500 ;
      RECT 0.7000 80.8500 461.8000 81.1500 ;
      RECT 0.0000 79.1500 461.8000 80.8500 ;
      RECT 0.7000 78.8500 461.8000 79.1500 ;
      RECT 0.0000 77.1500 461.8000 78.8500 ;
      RECT 0.7000 76.8500 461.8000 77.1500 ;
      RECT 0.0000 75.1500 461.8000 76.8500 ;
      RECT 0.7000 74.8500 461.8000 75.1500 ;
      RECT 0.0000 73.1500 461.8000 74.8500 ;
      RECT 0.7000 72.8500 461.8000 73.1500 ;
      RECT 0.0000 71.1500 461.8000 72.8500 ;
      RECT 0.7000 70.8500 461.8000 71.1500 ;
      RECT 0.0000 69.1500 461.8000 70.8500 ;
      RECT 0.7000 68.8500 461.8000 69.1500 ;
      RECT 0.0000 67.1500 461.8000 68.8500 ;
      RECT 0.7000 66.8500 461.8000 67.1500 ;
      RECT 0.0000 65.1500 461.8000 66.8500 ;
      RECT 0.7000 64.8500 461.8000 65.1500 ;
      RECT 0.0000 63.1500 461.8000 64.8500 ;
      RECT 0.7000 62.8500 461.8000 63.1500 ;
      RECT 0.0000 61.1500 461.8000 62.8500 ;
      RECT 0.7000 60.8500 461.8000 61.1500 ;
      RECT 0.0000 59.1500 461.8000 60.8500 ;
      RECT 0.7000 58.8500 461.8000 59.1500 ;
      RECT 0.0000 57.1500 461.8000 58.8500 ;
      RECT 0.7000 56.8500 461.8000 57.1500 ;
      RECT 0.0000 55.1500 461.8000 56.8500 ;
      RECT 0.7000 54.8500 461.8000 55.1500 ;
      RECT 0.0000 0.0000 461.8000 54.8500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 461.8000 459.2000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 461.8000 459.2000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 461.8000 459.2000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 461.8000 459.2000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 461.8000 459.2000 ;
  END
END fullchip

END LIBRARY
