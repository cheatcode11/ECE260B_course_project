// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// Please do not spread this code without permission 
module core (clk, sum_out, mem_in, out, inst, reset);

parameter col = 8;
parameter bw = 8;
parameter bw_psum = 2*bw+4;
parameter pr = 8;

output [bw_psum+3:0] sum_out;
output [bw_psum*col-1:0] out;
wire   [bw_psum*col-1:0] pmem_out;
input  [pr*bw-1:0] mem_in;
input  clk;
// Ajay: Bitwidth of inst increase by two to control sfp
input  [21:0] inst; 
input  reset;

wire  [pr*bw-1:0] mac_in;
wire  [pr*bw-1:0] kmem_out;
wire  [pr*bw-1:0] qmem_out;
wire  [bw_psum*col-1:0] pmem_in;
wire  [bw_psum*col-1:0] fifo_out;
// Output of SFP
wire  [bw_psum*col-1:0] sfp_out;
wire  [bw_psum*col-1:0] array_out;
wire  [bw_psum*col-1:0] fifo_sfp_out;  // New FIFO output between SFP and PMEM
wire  [col-1:0] fifo_wr;
wire  ofifo_rd;
wire [2:0] qkmem_add;
wire [2:0] pmem_add;

wire  qmem_rd;
wire  qmem_wr; 
wire  kmem_rd;
wire  kmem_wr; 
wire  pmem_rd;
wire  pmem_wr; 

assign ofifo_rd = inst[16];
assign qkmem_add = inst[15:12];
assign pmem_add = inst[11:8];

assign qmem_rd = inst[5];
assign qmem_wr = inst[4];
assign kmem_rd = inst[3];
assign kmem_wr = inst[2];
assign pmem_rd = inst[1];
assign pmem_wr = inst[0];

assign mac_in  = inst[6] ? kmem_out : qmem_out;
//assign pmem_in = fifo_sfp_out; // Now PMEM gets data from second FIFO

assign pmem_in = normalized_out; // Now PMEM gets data from second FIFO
// -----   SFP params -------
// Input of SFP
wire [bw_psum*col-1:0] to_normalize;
// Output of SFP
wire [bw_psum*col-1:0] normalized_out;
assign to_normalize = fifo_out;
assign out = pmem_out;
wire div = inst[17]; 
wire acc = inst[18];
wire [col-1:0] sfp_pmem_wr = inst[19];
wire fifo_ext_rd = 1'b0;
wire sum_in[24:0];
wire [23:0] sum_to_other_core; 

mac_array #(.bw(bw), .bw_psum(bw_psum), .col(col), .pr(pr)) mac_array_instance (
        .in(mac_in), 
        .clk(clk), 
        .reset(reset), 
        .inst(inst[7:6]),     
        .fifo_wr(fifo_wr),     
	.out(array_out)
);

ofifo #(.bw(bw_psum), .col(col))  ofifo_inst (
        .reset(reset),
        .clk(clk),
        .in(array_out),
        .wr(fifo_wr),
        .rd(ofifo_rd),
        .o_valid(fifo_valid),
        .out(fifo_out)
);

sfp_row #(.bw(bw), .bw_psum(bw_psum), .col(col)) sfp_instance(
	.clk(clk),
	.div(div),
	.acc(acc), 
	.fifo_ext_rd(fifo_ext_rd),   // 1'b0
	.sum_in(24'b1),   // 24'b0
	.sfp_in(to_normalize),
	.sfp_out(normalized_out),
	.sum_out(sum_to_other_core)	
);
/*
// Second FIFO: Stores SFP output before PMEM
ofifo #(.bw(bw_psum), .col(col))  sfp_fifo_inst (
        .reset(reset),
        .clk(clk),
        .in(normalized_out),
        .wr(sfp_pmem_wr), // Write when SFP processing is done
        .rd(ofifo_rd),    // Read when PMEM is ready
        .o_valid(fifo_valid),
        .out(fifo_sfp_out) // Output goes to PMEM
);
*/
sram_w16 #(.sram_bit(pr*bw)) qmem_instance (
        .CLK(clk),
        .D(mem_in),
        .Q(qmem_out),
        .CEN(!(qmem_rd||qmem_wr)),
        .WEN(!qmem_wr), 
        .A(qkmem_add)
);

sram_w16 #(.sram_bit(pr*bw)) kmem_instance (
        .CLK(clk),
        .D(mem_in),
        .Q(kmem_out),
        .CEN(!(kmem_rd||kmem_wr)),
        .WEN(!kmem_wr), 
        .A(qkmem_add)
);

sram_w16 #(.sram_bit(col*bw_psum)) psum_mem_instance (
        .CLK(clk),
        .D(pmem_in),
        .Q(pmem_out),
        .CEN(!(pmem_rd||pmem_wr)),
        .WEN(!pmem_wr),
        .A(pmem_add)
);

  //////////// For printing purpose ////////////
  always @(posedge clk) begin
      //if(pmem_wr)
         //$display("Memory write to PSUM mem add %x %x ", pmem_add, pmem_in); 
  end

endmodule
