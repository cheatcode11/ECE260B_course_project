// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// Please do not spread this code without permission 
module mac_array_gated_c (clk, reset, in, out, fifo_wr, inst, q_zero, ld_done, exec_done, out_wr);

parameter col = 8;
parameter bw = 8;
parameter bw_psum = 2*bw+6;
parameter pr = 8;

output [bw_psum*col-1:0] out;
input  [pr*bw-1:0] in;
input  clk, reset;
input  [1:0] inst; // [1]: execute, [0]: load 
input [pr-1:0] q_zero;
output [col-1:0] fifo_wr;
output ld_done;
output exec_done;
output out_wr;

wire   [col*bw_psum-1:0] psum;
wire   [2*(col+1)-1:0] inst_temp;
wire   [2*(col+1)*bw*pr-1:0] q_temp;
wire   [(col+1)*pr-1:0] q_zero_connector;
wire   [col-1:0] load_ready_wire;

genvar i;

//for (i=0; i < col ; i=i+1) begin
//  assign fifo_wr[i] = inst_temp[2*i+1] ;
//end

assign inst_temp[1:0]    = inst;
assign q_temp[bw*pr-1:0] = in;
assign q_zero_connector[pr-1:0] = q_zero;


for (i=1; i < col+1 ; i=i+1) begin : col_idx
   mac_col_gated_c #(.bw(bw), .bw_psum(bw_psum), .pr(pr), .col_id(i)) mac_col_inst (
        .q_in( q_temp[pr*bw*i-1    :pr*bw*(i-1)]), 
        .q_out(q_temp[pr*bw*(i+1)-1:pr*bw*i]), 
        .clk(clk), 
        .reset(reset), 
        .fifo_wr(fifo_wr[i-1]),
        .i_inst(inst_temp[2*i-1:2*(i-1)]),     
        .o_inst(inst_temp[2*(i+1)-1:2*(i)]),     
	.out(out[bw_psum*i-1 : bw_psum*(i-1)]),
	.q_zero(q_zero_connector[i*pr-1:(i-1)*pr]),
	.q_zero_out(q_zero_connector[(i+1)*pr-1:(i)*pr]),
	.load_ready(load_ready_wire[i-1])
   );
end 

assign ld_done = ~|load_ready_wire;
assign exec_done = (fifo_wr == 8'b00000111)? 1'b1: 1'b0;
assign out_wr = ~|fifo_wr;

endmodule

