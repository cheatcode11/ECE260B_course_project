##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sun Mar 16 01:34:20 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16
  CLASS BLOCK ;
  SIZE 678.6000 BY 53.8000 ;
  FOREIGN sram_w16 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.7500 0.8000 20.8500 ;
    END
  END CLK
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 593.0500 0.0000 593.1500 0.8000 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 589.0500 0.0000 589.1500 0.8000 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 585.0500 0.0000 585.1500 0.8000 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 581.0500 0.0000 581.1500 0.8000 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 577.0500 0.0000 577.1500 0.8000 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 573.0500 0.0000 573.1500 0.8000 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 569.0500 0.0000 569.1500 0.8000 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 565.0500 0.0000 565.1500 0.8000 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 561.0500 0.0000 561.1500 0.8000 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 557.0500 0.0000 557.1500 0.8000 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 553.0500 0.0000 553.1500 0.8000 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 549.0500 0.0000 549.1500 0.8000 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 545.0500 0.0000 545.1500 0.8000 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 541.0500 0.0000 541.1500 0.8000 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 537.0500 0.0000 537.1500 0.8000 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 533.0500 0.0000 533.1500 0.8000 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 529.0500 0.0000 529.1500 0.8000 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 525.0500 0.0000 525.1500 0.8000 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 521.0500 0.0000 521.1500 0.8000 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 517.0500 0.0000 517.1500 0.8000 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 513.0500 0.0000 513.1500 0.8000 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 509.0500 0.0000 509.1500 0.8000 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 505.0500 0.0000 505.1500 0.8000 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 501.0500 0.0000 501.1500 0.8000 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 497.0500 0.0000 497.1500 0.8000 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 493.0500 0.0000 493.1500 0.8000 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 489.0500 0.0000 489.1500 0.8000 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 485.0500 0.0000 485.1500 0.8000 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 481.0500 0.0000 481.1500 0.8000 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 477.0500 0.0000 477.1500 0.8000 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 473.0500 0.0000 473.1500 0.8000 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 469.0500 0.0000 469.1500 0.8000 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 465.0500 0.0000 465.1500 0.8000 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 461.0500 0.0000 461.1500 0.8000 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 457.0500 0.0000 457.1500 0.8000 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 453.0500 0.0000 453.1500 0.8000 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 449.0500 0.0000 449.1500 0.8000 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 445.0500 0.0000 445.1500 0.8000 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 441.0500 0.0000 441.1500 0.8000 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 437.0500 0.0000 437.1500 0.8000 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 433.0500 0.0000 433.1500 0.8000 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 429.0500 0.0000 429.1500 0.8000 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 425.0500 0.0000 425.1500 0.8000 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 421.0500 0.0000 421.1500 0.8000 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 417.0500 0.0000 417.1500 0.8000 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 413.0500 0.0000 413.1500 0.8000 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 409.0500 0.0000 409.1500 0.8000 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.0500 0.0000 405.1500 0.8000 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 401.0500 0.0000 401.1500 0.8000 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.0500 0.0000 397.1500 0.8000 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 393.0500 0.0000 393.1500 0.8000 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 389.0500 0.0000 389.1500 0.8000 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 385.0500 0.0000 385.1500 0.8000 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 381.0500 0.0000 381.1500 0.8000 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 377.0500 0.0000 377.1500 0.8000 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 373.0500 0.0000 373.1500 0.8000 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.0500 0.0000 369.1500 0.8000 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 365.0500 0.0000 365.1500 0.8000 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.0500 0.0000 361.1500 0.8000 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.0500 0.0000 357.1500 0.8000 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.0500 0.0000 353.1500 0.8000 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.0500 0.0000 349.1500 0.8000 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.0500 0.0000 345.1500 0.8000 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.0500 0.0000 341.1500 0.8000 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.0500 0.0000 337.1500 0.8000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.0500 0.0000 333.1500 0.8000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.0500 0.0000 329.1500 0.8000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.0500 0.0000 325.1500 0.8000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.0500 0.0000 321.1500 0.8000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.0500 0.0000 317.1500 0.8000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.0500 0.0000 313.1500 0.8000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.0500 0.0000 309.1500 0.8000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 305.0500 0.0000 305.1500 0.8000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 301.0500 0.0000 301.1500 0.8000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 297.0500 0.0000 297.1500 0.8000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 293.0500 0.0000 293.1500 0.8000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 289.0500 0.0000 289.1500 0.8000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 285.0500 0.0000 285.1500 0.8000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 281.0500 0.0000 281.1500 0.8000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.0500 0.0000 277.1500 0.8000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.0500 0.0000 273.1500 0.8000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 269.0500 0.0000 269.1500 0.8000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 265.0500 0.0000 265.1500 0.8000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 261.0500 0.0000 261.1500 0.8000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 257.0500 0.0000 257.1500 0.8000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 253.0500 0.0000 253.1500 0.8000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 249.0500 0.0000 249.1500 0.8000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 245.0500 0.0000 245.1500 0.8000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.0500 0.0000 241.1500 0.8000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.0500 0.0000 237.1500 0.8000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.0500 0.0000 233.1500 0.8000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 229.0500 0.0000 229.1500 0.8000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 225.0500 0.0000 225.1500 0.8000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 221.0500 0.0000 221.1500 0.8000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.0500 0.0000 217.1500 0.8000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.0500 0.0000 213.1500 0.8000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.0500 0.0000 209.1500 0.8000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.0500 0.0000 205.1500 0.8000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.0500 0.0000 201.1500 0.8000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.0500 0.0000 197.1500 0.8000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.0500 0.0000 193.1500 0.8000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.0500 0.0000 189.1500 0.8000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 185.0500 0.0000 185.1500 0.8000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.0500 0.0000 181.1500 0.8000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.0500 0.0000 177.1500 0.8000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.0500 0.0000 173.1500 0.8000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.0500 0.0000 169.1500 0.8000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.0500 0.0000 165.1500 0.8000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.0500 0.0000 161.1500 0.8000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.0500 0.0000 157.1500 0.8000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.0500 0.0000 153.1500 0.8000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.0500 0.0000 149.1500 0.8000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.0500 0.0000 145.1500 0.8000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.0500 0.0000 141.1500 0.8000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.0500 0.0000 137.1500 0.8000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.0500 0.0000 133.1500 0.8000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.0500 0.0000 129.1500 0.8000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.0500 0.0000 125.1500 0.8000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.0500 0.0000 121.1500 0.8000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.0500 0.0000 117.1500 0.8000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.0500 0.0000 113.1500 0.8000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.0500 0.0000 109.1500 0.8000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.0500 0.0000 105.1500 0.8000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.0500 0.0000 101.1500 0.8000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.0500 0.0000 97.1500 0.8000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.0500 0.0000 93.1500 0.8000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.0500 0.0000 89.1500 0.8000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.0500 0.0000 85.1500 0.8000 ;
    END
  END D[0]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 593.0500 53.0000 593.1500 53.8000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 589.0500 53.0000 589.1500 53.8000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 585.0500 53.0000 585.1500 53.8000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 581.0500 53.0000 581.1500 53.8000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 577.0500 53.0000 577.1500 53.8000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 573.0500 53.0000 573.1500 53.8000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 569.0500 53.0000 569.1500 53.8000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 565.0500 53.0000 565.1500 53.8000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 561.0500 53.0000 561.1500 53.8000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 557.0500 53.0000 557.1500 53.8000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 553.0500 53.0000 553.1500 53.8000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 549.0500 53.0000 549.1500 53.8000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 545.0500 53.0000 545.1500 53.8000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 541.0500 53.0000 541.1500 53.8000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 537.0500 53.0000 537.1500 53.8000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 533.0500 53.0000 533.1500 53.8000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 529.0500 53.0000 529.1500 53.8000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 525.0500 53.0000 525.1500 53.8000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 521.0500 53.0000 521.1500 53.8000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 517.0500 53.0000 517.1500 53.8000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 513.0500 53.0000 513.1500 53.8000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 509.0500 53.0000 509.1500 53.8000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 505.0500 53.0000 505.1500 53.8000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 501.0500 53.0000 501.1500 53.8000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 497.0500 53.0000 497.1500 53.8000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 493.0500 53.0000 493.1500 53.8000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 489.0500 53.0000 489.1500 53.8000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 485.0500 53.0000 485.1500 53.8000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 481.0500 53.0000 481.1500 53.8000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 477.0500 53.0000 477.1500 53.8000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 473.0500 53.0000 473.1500 53.8000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 469.0500 53.0000 469.1500 53.8000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 465.0500 53.0000 465.1500 53.8000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 461.0500 53.0000 461.1500 53.8000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 457.0500 53.0000 457.1500 53.8000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 453.0500 53.0000 453.1500 53.8000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 449.0500 53.0000 449.1500 53.8000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 445.0500 53.0000 445.1500 53.8000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 441.0500 53.0000 441.1500 53.8000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 437.0500 53.0000 437.1500 53.8000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 433.0500 53.0000 433.1500 53.8000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 429.0500 53.0000 429.1500 53.8000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 425.0500 53.0000 425.1500 53.8000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 421.0500 53.0000 421.1500 53.8000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 417.0500 53.0000 417.1500 53.8000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 413.0500 53.0000 413.1500 53.8000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 409.0500 53.0000 409.1500 53.8000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.0500 53.0000 405.1500 53.8000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 401.0500 53.0000 401.1500 53.8000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.0500 53.0000 397.1500 53.8000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 393.0500 53.0000 393.1500 53.8000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 389.0500 53.0000 389.1500 53.8000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 385.0500 53.0000 385.1500 53.8000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 381.0500 53.0000 381.1500 53.8000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 377.0500 53.0000 377.1500 53.8000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 373.0500 53.0000 373.1500 53.8000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.0500 53.0000 369.1500 53.8000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 365.0500 53.0000 365.1500 53.8000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.0500 53.0000 361.1500 53.8000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.0500 53.0000 357.1500 53.8000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.0500 53.0000 353.1500 53.8000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.0500 53.0000 349.1500 53.8000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.0500 53.0000 345.1500 53.8000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.0500 53.0000 341.1500 53.8000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.0500 53.0000 337.1500 53.8000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.0500 53.0000 333.1500 53.8000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.0500 53.0000 329.1500 53.8000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.0500 53.0000 325.1500 53.8000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.0500 53.0000 321.1500 53.8000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.0500 53.0000 317.1500 53.8000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 313.0500 53.0000 313.1500 53.8000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.0500 53.0000 309.1500 53.8000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 305.0500 53.0000 305.1500 53.8000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 301.0500 53.0000 301.1500 53.8000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 297.0500 53.0000 297.1500 53.8000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 293.0500 53.0000 293.1500 53.8000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 289.0500 53.0000 289.1500 53.8000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 285.0500 53.0000 285.1500 53.8000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 281.0500 53.0000 281.1500 53.8000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.0500 53.0000 277.1500 53.8000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.0500 53.0000 273.1500 53.8000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 269.0500 53.0000 269.1500 53.8000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 265.0500 53.0000 265.1500 53.8000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 261.0500 53.0000 261.1500 53.8000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 257.0500 53.0000 257.1500 53.8000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 253.0500 53.0000 253.1500 53.8000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 249.0500 53.0000 249.1500 53.8000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 245.0500 53.0000 245.1500 53.8000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.0500 53.0000 241.1500 53.8000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.0500 53.0000 237.1500 53.8000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.0500 53.0000 233.1500 53.8000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 229.0500 53.0000 229.1500 53.8000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 225.0500 53.0000 225.1500 53.8000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 221.0500 53.0000 221.1500 53.8000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.0500 53.0000 217.1500 53.8000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.0500 53.0000 213.1500 53.8000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.0500 53.0000 209.1500 53.8000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.0500 53.0000 205.1500 53.8000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.0500 53.0000 201.1500 53.8000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.0500 53.0000 197.1500 53.8000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.0500 53.0000 193.1500 53.8000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.0500 53.0000 189.1500 53.8000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 185.0500 53.0000 185.1500 53.8000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.0500 53.0000 181.1500 53.8000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.0500 53.0000 177.1500 53.8000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.0500 53.0000 173.1500 53.8000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.0500 53.0000 169.1500 53.8000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.0500 53.0000 165.1500 53.8000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.0500 53.0000 161.1500 53.8000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.0500 53.0000 157.1500 53.8000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.0500 53.0000 153.1500 53.8000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.0500 53.0000 149.1500 53.8000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.0500 53.0000 145.1500 53.8000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.0500 53.0000 141.1500 53.8000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.0500 53.0000 137.1500 53.8000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.0500 53.0000 133.1500 53.8000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.0500 53.0000 129.1500 53.8000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.0500 53.0000 125.1500 53.8000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.0500 53.0000 121.1500 53.8000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.0500 53.0000 117.1500 53.8000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.0500 53.0000 113.1500 53.8000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.0500 53.0000 109.1500 53.8000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.0500 53.0000 105.1500 53.8000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.0500 53.0000 101.1500 53.8000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.0500 53.0000 97.1500 53.8000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.0500 53.0000 93.1500 53.8000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.0500 53.0000 89.1500 53.8000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.0500 53.0000 85.1500 53.8000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.7500 0.8000 16.8500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 36.7500 0.8000 36.8500 ;
    END
  END WEN
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.7500 0.8000 32.8500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.7500 0.8000 28.8500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.7500 0.8000 24.8500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 20.0000 8.0000 21.0000 45.8000 ;
        RECT 88.5550 8.0000 89.5550 45.8000 ;
        RECT 157.1100 8.0000 158.1100 45.8000 ;
        RECT 225.6650 8.0000 226.6650 45.8000 ;
        RECT 294.2200 8.0000 295.2200 45.8000 ;
        RECT 362.7750 8.0000 363.7750 45.8000 ;
        RECT 431.3300 8.0000 432.3300 45.8000 ;
        RECT 499.8850 8.0000 500.8850 45.8000 ;
        RECT 568.4400 8.0000 569.4400 45.8000 ;
        RECT 636.9950 8.0000 637.9950 45.8000 ;
        RECT 20.0000 45.6350 21.0000 45.9650 ;
        RECT 88.5550 45.6350 89.5550 45.9650 ;
        RECT 157.1100 45.6350 158.1100 45.9650 ;
        RECT 225.6650 45.6350 226.6650 45.9650 ;
        RECT 294.2200 45.6350 295.2200 45.9650 ;
        RECT 362.7750 45.6350 363.7750 45.9650 ;
        RECT 431.3300 45.6350 432.3300 45.9650 ;
        RECT 499.8850 45.6350 500.8850 45.9650 ;
        RECT 568.4400 45.6350 569.4400 45.9650 ;
        RECT 636.9950 45.6350 637.9950 45.9650 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 22.0000 8.0000 23.0000 45.8000 ;
        RECT 90.5550 8.0000 91.5550 45.8000 ;
        RECT 159.1100 8.0000 160.1100 45.8000 ;
        RECT 227.6650 8.0000 228.6650 45.8000 ;
        RECT 296.2200 8.0000 297.2200 45.8000 ;
        RECT 364.7750 8.0000 365.7750 45.8000 ;
        RECT 433.3300 8.0000 434.3300 45.8000 ;
        RECT 501.8850 8.0000 502.8850 45.8000 ;
        RECT 570.4400 8.0000 571.4400 45.8000 ;
        RECT 638.9950 8.0000 639.9950 45.8000 ;
        RECT 22.0000 7.8350 23.0000 8.1650 ;
        RECT 90.5550 7.8350 91.5550 8.1650 ;
        RECT 159.1100 7.8350 160.1100 8.1650 ;
        RECT 227.6650 7.8350 228.6650 8.1650 ;
        RECT 296.2200 7.8350 297.2200 8.1650 ;
        RECT 364.7750 7.8350 365.7750 8.1650 ;
        RECT 433.3300 7.8350 434.3300 8.1650 ;
        RECT 501.8850 7.8350 502.8850 8.1650 ;
        RECT 570.4400 7.8350 571.4400 8.1650 ;
        RECT 638.9950 7.8350 639.9950 8.1650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 678.6000 53.8000 ;
    LAYER M2 ;
      RECT 593.2500 52.9000 678.6000 53.8000 ;
      RECT 589.2500 52.9000 592.9500 53.8000 ;
      RECT 585.2500 52.9000 588.9500 53.8000 ;
      RECT 581.2500 52.9000 584.9500 53.8000 ;
      RECT 577.2500 52.9000 580.9500 53.8000 ;
      RECT 573.2500 52.9000 576.9500 53.8000 ;
      RECT 569.2500 52.9000 572.9500 53.8000 ;
      RECT 565.2500 52.9000 568.9500 53.8000 ;
      RECT 561.2500 52.9000 564.9500 53.8000 ;
      RECT 557.2500 52.9000 560.9500 53.8000 ;
      RECT 553.2500 52.9000 556.9500 53.8000 ;
      RECT 549.2500 52.9000 552.9500 53.8000 ;
      RECT 545.2500 52.9000 548.9500 53.8000 ;
      RECT 541.2500 52.9000 544.9500 53.8000 ;
      RECT 537.2500 52.9000 540.9500 53.8000 ;
      RECT 533.2500 52.9000 536.9500 53.8000 ;
      RECT 529.2500 52.9000 532.9500 53.8000 ;
      RECT 525.2500 52.9000 528.9500 53.8000 ;
      RECT 521.2500 52.9000 524.9500 53.8000 ;
      RECT 517.2500 52.9000 520.9500 53.8000 ;
      RECT 513.2500 52.9000 516.9500 53.8000 ;
      RECT 509.2500 52.9000 512.9500 53.8000 ;
      RECT 505.2500 52.9000 508.9500 53.8000 ;
      RECT 501.2500 52.9000 504.9500 53.8000 ;
      RECT 497.2500 52.9000 500.9500 53.8000 ;
      RECT 493.2500 52.9000 496.9500 53.8000 ;
      RECT 489.2500 52.9000 492.9500 53.8000 ;
      RECT 485.2500 52.9000 488.9500 53.8000 ;
      RECT 481.2500 52.9000 484.9500 53.8000 ;
      RECT 477.2500 52.9000 480.9500 53.8000 ;
      RECT 473.2500 52.9000 476.9500 53.8000 ;
      RECT 469.2500 52.9000 472.9500 53.8000 ;
      RECT 465.2500 52.9000 468.9500 53.8000 ;
      RECT 461.2500 52.9000 464.9500 53.8000 ;
      RECT 457.2500 52.9000 460.9500 53.8000 ;
      RECT 453.2500 52.9000 456.9500 53.8000 ;
      RECT 449.2500 52.9000 452.9500 53.8000 ;
      RECT 445.2500 52.9000 448.9500 53.8000 ;
      RECT 441.2500 52.9000 444.9500 53.8000 ;
      RECT 437.2500 52.9000 440.9500 53.8000 ;
      RECT 433.2500 52.9000 436.9500 53.8000 ;
      RECT 429.2500 52.9000 432.9500 53.8000 ;
      RECT 425.2500 52.9000 428.9500 53.8000 ;
      RECT 421.2500 52.9000 424.9500 53.8000 ;
      RECT 417.2500 52.9000 420.9500 53.8000 ;
      RECT 413.2500 52.9000 416.9500 53.8000 ;
      RECT 409.2500 52.9000 412.9500 53.8000 ;
      RECT 405.2500 52.9000 408.9500 53.8000 ;
      RECT 401.2500 52.9000 404.9500 53.8000 ;
      RECT 397.2500 52.9000 400.9500 53.8000 ;
      RECT 393.2500 52.9000 396.9500 53.8000 ;
      RECT 389.2500 52.9000 392.9500 53.8000 ;
      RECT 385.2500 52.9000 388.9500 53.8000 ;
      RECT 381.2500 52.9000 384.9500 53.8000 ;
      RECT 377.2500 52.9000 380.9500 53.8000 ;
      RECT 373.2500 52.9000 376.9500 53.8000 ;
      RECT 369.2500 52.9000 372.9500 53.8000 ;
      RECT 365.2500 52.9000 368.9500 53.8000 ;
      RECT 361.2500 52.9000 364.9500 53.8000 ;
      RECT 357.2500 52.9000 360.9500 53.8000 ;
      RECT 353.2500 52.9000 356.9500 53.8000 ;
      RECT 349.2500 52.9000 352.9500 53.8000 ;
      RECT 345.2500 52.9000 348.9500 53.8000 ;
      RECT 341.2500 52.9000 344.9500 53.8000 ;
      RECT 337.2500 52.9000 340.9500 53.8000 ;
      RECT 333.2500 52.9000 336.9500 53.8000 ;
      RECT 329.2500 52.9000 332.9500 53.8000 ;
      RECT 325.2500 52.9000 328.9500 53.8000 ;
      RECT 321.2500 52.9000 324.9500 53.8000 ;
      RECT 317.2500 52.9000 320.9500 53.8000 ;
      RECT 313.2500 52.9000 316.9500 53.8000 ;
      RECT 309.2500 52.9000 312.9500 53.8000 ;
      RECT 305.2500 52.9000 308.9500 53.8000 ;
      RECT 301.2500 52.9000 304.9500 53.8000 ;
      RECT 297.2500 52.9000 300.9500 53.8000 ;
      RECT 293.2500 52.9000 296.9500 53.8000 ;
      RECT 289.2500 52.9000 292.9500 53.8000 ;
      RECT 285.2500 52.9000 288.9500 53.8000 ;
      RECT 281.2500 52.9000 284.9500 53.8000 ;
      RECT 277.2500 52.9000 280.9500 53.8000 ;
      RECT 273.2500 52.9000 276.9500 53.8000 ;
      RECT 269.2500 52.9000 272.9500 53.8000 ;
      RECT 265.2500 52.9000 268.9500 53.8000 ;
      RECT 261.2500 52.9000 264.9500 53.8000 ;
      RECT 257.2500 52.9000 260.9500 53.8000 ;
      RECT 253.2500 52.9000 256.9500 53.8000 ;
      RECT 249.2500 52.9000 252.9500 53.8000 ;
      RECT 245.2500 52.9000 248.9500 53.8000 ;
      RECT 241.2500 52.9000 244.9500 53.8000 ;
      RECT 237.2500 52.9000 240.9500 53.8000 ;
      RECT 233.2500 52.9000 236.9500 53.8000 ;
      RECT 229.2500 52.9000 232.9500 53.8000 ;
      RECT 225.2500 52.9000 228.9500 53.8000 ;
      RECT 221.2500 52.9000 224.9500 53.8000 ;
      RECT 217.2500 52.9000 220.9500 53.8000 ;
      RECT 213.2500 52.9000 216.9500 53.8000 ;
      RECT 209.2500 52.9000 212.9500 53.8000 ;
      RECT 205.2500 52.9000 208.9500 53.8000 ;
      RECT 201.2500 52.9000 204.9500 53.8000 ;
      RECT 197.2500 52.9000 200.9500 53.8000 ;
      RECT 193.2500 52.9000 196.9500 53.8000 ;
      RECT 189.2500 52.9000 192.9500 53.8000 ;
      RECT 185.2500 52.9000 188.9500 53.8000 ;
      RECT 181.2500 52.9000 184.9500 53.8000 ;
      RECT 177.2500 52.9000 180.9500 53.8000 ;
      RECT 173.2500 52.9000 176.9500 53.8000 ;
      RECT 169.2500 52.9000 172.9500 53.8000 ;
      RECT 165.2500 52.9000 168.9500 53.8000 ;
      RECT 161.2500 52.9000 164.9500 53.8000 ;
      RECT 157.2500 52.9000 160.9500 53.8000 ;
      RECT 153.2500 52.9000 156.9500 53.8000 ;
      RECT 149.2500 52.9000 152.9500 53.8000 ;
      RECT 145.2500 52.9000 148.9500 53.8000 ;
      RECT 141.2500 52.9000 144.9500 53.8000 ;
      RECT 137.2500 52.9000 140.9500 53.8000 ;
      RECT 133.2500 52.9000 136.9500 53.8000 ;
      RECT 129.2500 52.9000 132.9500 53.8000 ;
      RECT 125.2500 52.9000 128.9500 53.8000 ;
      RECT 121.2500 52.9000 124.9500 53.8000 ;
      RECT 117.2500 52.9000 120.9500 53.8000 ;
      RECT 113.2500 52.9000 116.9500 53.8000 ;
      RECT 109.2500 52.9000 112.9500 53.8000 ;
      RECT 105.2500 52.9000 108.9500 53.8000 ;
      RECT 101.2500 52.9000 104.9500 53.8000 ;
      RECT 97.2500 52.9000 100.9500 53.8000 ;
      RECT 93.2500 52.9000 96.9500 53.8000 ;
      RECT 89.2500 52.9000 92.9500 53.8000 ;
      RECT 85.2500 52.9000 88.9500 53.8000 ;
      RECT 0.0000 52.9000 84.9500 53.8000 ;
      RECT 0.0000 0.9000 678.6000 52.9000 ;
      RECT 593.2500 0.0000 678.6000 0.9000 ;
      RECT 589.2500 0.0000 592.9500 0.9000 ;
      RECT 585.2500 0.0000 588.9500 0.9000 ;
      RECT 581.2500 0.0000 584.9500 0.9000 ;
      RECT 577.2500 0.0000 580.9500 0.9000 ;
      RECT 573.2500 0.0000 576.9500 0.9000 ;
      RECT 569.2500 0.0000 572.9500 0.9000 ;
      RECT 565.2500 0.0000 568.9500 0.9000 ;
      RECT 561.2500 0.0000 564.9500 0.9000 ;
      RECT 557.2500 0.0000 560.9500 0.9000 ;
      RECT 553.2500 0.0000 556.9500 0.9000 ;
      RECT 549.2500 0.0000 552.9500 0.9000 ;
      RECT 545.2500 0.0000 548.9500 0.9000 ;
      RECT 541.2500 0.0000 544.9500 0.9000 ;
      RECT 537.2500 0.0000 540.9500 0.9000 ;
      RECT 533.2500 0.0000 536.9500 0.9000 ;
      RECT 529.2500 0.0000 532.9500 0.9000 ;
      RECT 525.2500 0.0000 528.9500 0.9000 ;
      RECT 521.2500 0.0000 524.9500 0.9000 ;
      RECT 517.2500 0.0000 520.9500 0.9000 ;
      RECT 513.2500 0.0000 516.9500 0.9000 ;
      RECT 509.2500 0.0000 512.9500 0.9000 ;
      RECT 505.2500 0.0000 508.9500 0.9000 ;
      RECT 501.2500 0.0000 504.9500 0.9000 ;
      RECT 497.2500 0.0000 500.9500 0.9000 ;
      RECT 493.2500 0.0000 496.9500 0.9000 ;
      RECT 489.2500 0.0000 492.9500 0.9000 ;
      RECT 485.2500 0.0000 488.9500 0.9000 ;
      RECT 481.2500 0.0000 484.9500 0.9000 ;
      RECT 477.2500 0.0000 480.9500 0.9000 ;
      RECT 473.2500 0.0000 476.9500 0.9000 ;
      RECT 469.2500 0.0000 472.9500 0.9000 ;
      RECT 465.2500 0.0000 468.9500 0.9000 ;
      RECT 461.2500 0.0000 464.9500 0.9000 ;
      RECT 457.2500 0.0000 460.9500 0.9000 ;
      RECT 453.2500 0.0000 456.9500 0.9000 ;
      RECT 449.2500 0.0000 452.9500 0.9000 ;
      RECT 445.2500 0.0000 448.9500 0.9000 ;
      RECT 441.2500 0.0000 444.9500 0.9000 ;
      RECT 437.2500 0.0000 440.9500 0.9000 ;
      RECT 433.2500 0.0000 436.9500 0.9000 ;
      RECT 429.2500 0.0000 432.9500 0.9000 ;
      RECT 425.2500 0.0000 428.9500 0.9000 ;
      RECT 421.2500 0.0000 424.9500 0.9000 ;
      RECT 417.2500 0.0000 420.9500 0.9000 ;
      RECT 413.2500 0.0000 416.9500 0.9000 ;
      RECT 409.2500 0.0000 412.9500 0.9000 ;
      RECT 405.2500 0.0000 408.9500 0.9000 ;
      RECT 401.2500 0.0000 404.9500 0.9000 ;
      RECT 397.2500 0.0000 400.9500 0.9000 ;
      RECT 393.2500 0.0000 396.9500 0.9000 ;
      RECT 389.2500 0.0000 392.9500 0.9000 ;
      RECT 385.2500 0.0000 388.9500 0.9000 ;
      RECT 381.2500 0.0000 384.9500 0.9000 ;
      RECT 377.2500 0.0000 380.9500 0.9000 ;
      RECT 373.2500 0.0000 376.9500 0.9000 ;
      RECT 369.2500 0.0000 372.9500 0.9000 ;
      RECT 365.2500 0.0000 368.9500 0.9000 ;
      RECT 361.2500 0.0000 364.9500 0.9000 ;
      RECT 357.2500 0.0000 360.9500 0.9000 ;
      RECT 353.2500 0.0000 356.9500 0.9000 ;
      RECT 349.2500 0.0000 352.9500 0.9000 ;
      RECT 345.2500 0.0000 348.9500 0.9000 ;
      RECT 341.2500 0.0000 344.9500 0.9000 ;
      RECT 337.2500 0.0000 340.9500 0.9000 ;
      RECT 333.2500 0.0000 336.9500 0.9000 ;
      RECT 329.2500 0.0000 332.9500 0.9000 ;
      RECT 325.2500 0.0000 328.9500 0.9000 ;
      RECT 321.2500 0.0000 324.9500 0.9000 ;
      RECT 317.2500 0.0000 320.9500 0.9000 ;
      RECT 313.2500 0.0000 316.9500 0.9000 ;
      RECT 309.2500 0.0000 312.9500 0.9000 ;
      RECT 305.2500 0.0000 308.9500 0.9000 ;
      RECT 301.2500 0.0000 304.9500 0.9000 ;
      RECT 297.2500 0.0000 300.9500 0.9000 ;
      RECT 293.2500 0.0000 296.9500 0.9000 ;
      RECT 289.2500 0.0000 292.9500 0.9000 ;
      RECT 285.2500 0.0000 288.9500 0.9000 ;
      RECT 281.2500 0.0000 284.9500 0.9000 ;
      RECT 277.2500 0.0000 280.9500 0.9000 ;
      RECT 273.2500 0.0000 276.9500 0.9000 ;
      RECT 269.2500 0.0000 272.9500 0.9000 ;
      RECT 265.2500 0.0000 268.9500 0.9000 ;
      RECT 261.2500 0.0000 264.9500 0.9000 ;
      RECT 257.2500 0.0000 260.9500 0.9000 ;
      RECT 253.2500 0.0000 256.9500 0.9000 ;
      RECT 249.2500 0.0000 252.9500 0.9000 ;
      RECT 245.2500 0.0000 248.9500 0.9000 ;
      RECT 241.2500 0.0000 244.9500 0.9000 ;
      RECT 237.2500 0.0000 240.9500 0.9000 ;
      RECT 233.2500 0.0000 236.9500 0.9000 ;
      RECT 229.2500 0.0000 232.9500 0.9000 ;
      RECT 225.2500 0.0000 228.9500 0.9000 ;
      RECT 221.2500 0.0000 224.9500 0.9000 ;
      RECT 217.2500 0.0000 220.9500 0.9000 ;
      RECT 213.2500 0.0000 216.9500 0.9000 ;
      RECT 209.2500 0.0000 212.9500 0.9000 ;
      RECT 205.2500 0.0000 208.9500 0.9000 ;
      RECT 201.2500 0.0000 204.9500 0.9000 ;
      RECT 197.2500 0.0000 200.9500 0.9000 ;
      RECT 193.2500 0.0000 196.9500 0.9000 ;
      RECT 189.2500 0.0000 192.9500 0.9000 ;
      RECT 185.2500 0.0000 188.9500 0.9000 ;
      RECT 181.2500 0.0000 184.9500 0.9000 ;
      RECT 177.2500 0.0000 180.9500 0.9000 ;
      RECT 173.2500 0.0000 176.9500 0.9000 ;
      RECT 169.2500 0.0000 172.9500 0.9000 ;
      RECT 165.2500 0.0000 168.9500 0.9000 ;
      RECT 161.2500 0.0000 164.9500 0.9000 ;
      RECT 157.2500 0.0000 160.9500 0.9000 ;
      RECT 153.2500 0.0000 156.9500 0.9000 ;
      RECT 149.2500 0.0000 152.9500 0.9000 ;
      RECT 145.2500 0.0000 148.9500 0.9000 ;
      RECT 141.2500 0.0000 144.9500 0.9000 ;
      RECT 137.2500 0.0000 140.9500 0.9000 ;
      RECT 133.2500 0.0000 136.9500 0.9000 ;
      RECT 129.2500 0.0000 132.9500 0.9000 ;
      RECT 125.2500 0.0000 128.9500 0.9000 ;
      RECT 121.2500 0.0000 124.9500 0.9000 ;
      RECT 117.2500 0.0000 120.9500 0.9000 ;
      RECT 113.2500 0.0000 116.9500 0.9000 ;
      RECT 109.2500 0.0000 112.9500 0.9000 ;
      RECT 105.2500 0.0000 108.9500 0.9000 ;
      RECT 101.2500 0.0000 104.9500 0.9000 ;
      RECT 97.2500 0.0000 100.9500 0.9000 ;
      RECT 93.2500 0.0000 96.9500 0.9000 ;
      RECT 89.2500 0.0000 92.9500 0.9000 ;
      RECT 85.2500 0.0000 88.9500 0.9000 ;
      RECT 0.0000 0.0000 84.9500 0.9000 ;
    LAYER M3 ;
      RECT 0.0000 36.9500 678.6000 53.8000 ;
      RECT 0.9000 36.6500 678.6000 36.9500 ;
      RECT 0.0000 32.9500 678.6000 36.6500 ;
      RECT 0.9000 32.6500 678.6000 32.9500 ;
      RECT 0.0000 28.9500 678.6000 32.6500 ;
      RECT 0.9000 28.6500 678.6000 28.9500 ;
      RECT 0.0000 24.9500 678.6000 28.6500 ;
      RECT 0.9000 24.6500 678.6000 24.9500 ;
      RECT 0.0000 20.9500 678.6000 24.6500 ;
      RECT 0.9000 20.6500 678.6000 20.9500 ;
      RECT 0.0000 16.9500 678.6000 20.6500 ;
      RECT 0.9000 16.6500 678.6000 16.9500 ;
      RECT 0.0000 0.0000 678.6000 16.6500 ;
    LAYER M4 ;
      RECT 0.0000 46.1250 678.6000 53.8000 ;
      RECT 638.1550 45.9600 678.6000 46.1250 ;
      RECT 569.6000 45.9600 636.8350 46.1250 ;
      RECT 501.0450 45.9600 568.2800 46.1250 ;
      RECT 432.4900 45.9600 499.7250 46.1250 ;
      RECT 363.9350 45.9600 431.1700 46.1250 ;
      RECT 295.3800 45.9600 362.6150 46.1250 ;
      RECT 226.8250 45.9600 294.0600 46.1250 ;
      RECT 158.2700 45.9600 225.5050 46.1250 ;
      RECT 89.7150 45.9600 156.9500 46.1250 ;
      RECT 21.1600 45.9600 88.3950 46.1250 ;
      RECT 638.1550 7.8400 638.8350 45.9600 ;
      RECT 571.6000 7.8400 636.8350 45.9600 ;
      RECT 569.6000 7.8400 570.2800 45.9600 ;
      RECT 503.0450 7.8400 568.2800 45.9600 ;
      RECT 501.0450 7.8400 501.7250 45.9600 ;
      RECT 434.4900 7.8400 499.7250 45.9600 ;
      RECT 432.4900 7.8400 433.1700 45.9600 ;
      RECT 365.9350 7.8400 431.1700 45.9600 ;
      RECT 363.9350 7.8400 364.6150 45.9600 ;
      RECT 297.3800 7.8400 362.6150 45.9600 ;
      RECT 295.3800 7.8400 296.0600 45.9600 ;
      RECT 228.8250 7.8400 294.0600 45.9600 ;
      RECT 226.8250 7.8400 227.5050 45.9600 ;
      RECT 160.2700 7.8400 225.5050 45.9600 ;
      RECT 158.2700 7.8400 158.9500 45.9600 ;
      RECT 91.7150 7.8400 156.9500 45.9600 ;
      RECT 89.7150 7.8400 90.3950 45.9600 ;
      RECT 23.1600 7.8400 88.3950 45.9600 ;
      RECT 21.1600 7.8400 21.8400 45.9600 ;
      RECT 0.0000 7.8400 19.8400 46.1250 ;
      RECT 640.1550 7.6750 678.6000 45.9600 ;
      RECT 571.6000 7.6750 638.8350 7.8400 ;
      RECT 503.0450 7.6750 570.2800 7.8400 ;
      RECT 434.4900 7.6750 501.7250 7.8400 ;
      RECT 365.9350 7.6750 433.1700 7.8400 ;
      RECT 297.3800 7.6750 364.6150 7.8400 ;
      RECT 228.8250 7.6750 296.0600 7.8400 ;
      RECT 160.2700 7.6750 227.5050 7.8400 ;
      RECT 91.7150 7.6750 158.9500 7.8400 ;
      RECT 23.1600 7.6750 90.3950 7.8400 ;
      RECT 0.0000 7.6750 21.8400 7.8400 ;
      RECT 0.0000 0.0000 678.6000 7.6750 ;
  END
END sram_w16

END LIBRARY
