##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar 21 03:39:39 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16_2
  CLASS BLOCK ;
  SIZE 739.0000 BY 59.2000 ;
  FOREIGN sram_w16_2 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.3500 0.8000 23.4500 ;
    END
  END CLK
  PIN D[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 687.2500 0.0000 687.3500 0.8000 ;
    END
  END D[159]
  PIN D[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 683.2500 0.0000 683.3500 0.8000 ;
    END
  END D[158]
  PIN D[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 679.2500 0.0000 679.3500 0.8000 ;
    END
  END D[157]
  PIN D[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 675.2500 0.0000 675.3500 0.8000 ;
    END
  END D[156]
  PIN D[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 671.2500 0.0000 671.3500 0.8000 ;
    END
  END D[155]
  PIN D[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 667.2500 0.0000 667.3500 0.8000 ;
    END
  END D[154]
  PIN D[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 663.2500 0.0000 663.3500 0.8000 ;
    END
  END D[153]
  PIN D[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 659.2500 0.0000 659.3500 0.8000 ;
    END
  END D[152]
  PIN D[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 655.2500 0.0000 655.3500 0.8000 ;
    END
  END D[151]
  PIN D[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 651.2500 0.0000 651.3500 0.8000 ;
    END
  END D[150]
  PIN D[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 647.2500 0.0000 647.3500 0.8000 ;
    END
  END D[149]
  PIN D[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 643.2500 0.0000 643.3500 0.8000 ;
    END
  END D[148]
  PIN D[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 639.2500 0.0000 639.3500 0.8000 ;
    END
  END D[147]
  PIN D[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 635.2500 0.0000 635.3500 0.8000 ;
    END
  END D[146]
  PIN D[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 631.2500 0.0000 631.3500 0.8000 ;
    END
  END D[145]
  PIN D[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 627.2500 0.0000 627.3500 0.8000 ;
    END
  END D[144]
  PIN D[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 623.2500 0.0000 623.3500 0.8000 ;
    END
  END D[143]
  PIN D[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 619.2500 0.0000 619.3500 0.8000 ;
    END
  END D[142]
  PIN D[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 615.2500 0.0000 615.3500 0.8000 ;
    END
  END D[141]
  PIN D[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 611.2500 0.0000 611.3500 0.8000 ;
    END
  END D[140]
  PIN D[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 607.2500 0.0000 607.3500 0.8000 ;
    END
  END D[139]
  PIN D[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 603.2500 0.0000 603.3500 0.8000 ;
    END
  END D[138]
  PIN D[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 599.2500 0.0000 599.3500 0.8000 ;
    END
  END D[137]
  PIN D[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 595.2500 0.0000 595.3500 0.8000 ;
    END
  END D[136]
  PIN D[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 591.2500 0.0000 591.3500 0.8000 ;
    END
  END D[135]
  PIN D[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 587.2500 0.0000 587.3500 0.8000 ;
    END
  END D[134]
  PIN D[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 583.2500 0.0000 583.3500 0.8000 ;
    END
  END D[133]
  PIN D[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 579.2500 0.0000 579.3500 0.8000 ;
    END
  END D[132]
  PIN D[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 575.2500 0.0000 575.3500 0.8000 ;
    END
  END D[131]
  PIN D[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 571.2500 0.0000 571.3500 0.8000 ;
    END
  END D[130]
  PIN D[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 567.2500 0.0000 567.3500 0.8000 ;
    END
  END D[129]
  PIN D[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 563.2500 0.0000 563.3500 0.8000 ;
    END
  END D[128]
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 559.2500 0.0000 559.3500 0.8000 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 555.2500 0.0000 555.3500 0.8000 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 551.2500 0.0000 551.3500 0.8000 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 547.2500 0.0000 547.3500 0.8000 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 543.2500 0.0000 543.3500 0.8000 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 539.2500 0.0000 539.3500 0.8000 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 535.2500 0.0000 535.3500 0.8000 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 531.2500 0.0000 531.3500 0.8000 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 527.2500 0.0000 527.3500 0.8000 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 523.2500 0.0000 523.3500 0.8000 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 519.2500 0.0000 519.3500 0.8000 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 515.2500 0.0000 515.3500 0.8000 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 511.2500 0.0000 511.3500 0.8000 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 507.2500 0.0000 507.3500 0.8000 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 503.2500 0.0000 503.3500 0.8000 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 499.2500 0.0000 499.3500 0.8000 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 495.2500 0.0000 495.3500 0.8000 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 491.2500 0.0000 491.3500 0.8000 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 487.2500 0.0000 487.3500 0.8000 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 483.2500 0.0000 483.3500 0.8000 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 479.2500 0.0000 479.3500 0.8000 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 475.2500 0.0000 475.3500 0.8000 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 471.2500 0.0000 471.3500 0.8000 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 467.2500 0.0000 467.3500 0.8000 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 463.2500 0.0000 463.3500 0.8000 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 459.2500 0.0000 459.3500 0.8000 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 455.2500 0.0000 455.3500 0.8000 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 451.2500 0.0000 451.3500 0.8000 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.2500 0.0000 447.3500 0.8000 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.2500 0.0000 443.3500 0.8000 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.2500 0.0000 439.3500 0.8000 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.2500 0.0000 435.3500 0.8000 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 431.2500 0.0000 431.3500 0.8000 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.2500 0.0000 427.3500 0.8000 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.2500 0.0000 423.3500 0.8000 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.2500 0.0000 419.3500 0.8000 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.2500 0.0000 415.3500 0.8000 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 411.2500 0.0000 411.3500 0.8000 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.2500 0.0000 407.3500 0.8000 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.2500 0.0000 403.3500 0.8000 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.2500 0.0000 399.3500 0.8000 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.2500 0.0000 395.3500 0.8000 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.2500 0.0000 391.3500 0.8000 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.2500 0.0000 387.3500 0.8000 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.2500 0.0000 383.3500 0.8000 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 379.2500 0.0000 379.3500 0.8000 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.2500 0.0000 375.3500 0.8000 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.2500 0.0000 371.3500 0.8000 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.2500 0.0000 367.3500 0.8000 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.2500 0.0000 363.3500 0.8000 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.2500 0.0000 359.3500 0.8000 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.2500 0.0000 355.3500 0.8000 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.2500 0.0000 351.3500 0.8000 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.2500 0.0000 347.3500 0.8000 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.2500 0.0000 343.3500 0.8000 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.2500 0.0000 339.3500 0.8000 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.2500 0.0000 335.3500 0.8000 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.2500 0.0000 331.3500 0.8000 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.2500 0.0000 327.3500 0.8000 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.2500 0.0000 323.3500 0.8000 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.2500 0.0000 319.3500 0.8000 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.2500 0.0000 315.3500 0.8000 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.2500 0.0000 311.3500 0.8000 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.2500 0.0000 307.3500 0.8000 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.2500 0.0000 303.3500 0.8000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 299.2500 0.0000 299.3500 0.8000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.2500 0.0000 295.3500 0.8000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.2500 0.0000 291.3500 0.8000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 287.2500 0.0000 287.3500 0.8000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 283.2500 0.0000 283.3500 0.8000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 279.2500 0.0000 279.3500 0.8000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 275.2500 0.0000 275.3500 0.8000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 271.2500 0.0000 271.3500 0.8000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.2500 0.0000 267.3500 0.8000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 263.2500 0.0000 263.3500 0.8000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.2500 0.0000 259.3500 0.8000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.2500 0.0000 255.3500 0.8000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 251.2500 0.0000 251.3500 0.8000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.2500 0.0000 247.3500 0.8000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.2500 0.0000 243.3500 0.8000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 239.2500 0.0000 239.3500 0.8000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.2500 0.0000 235.3500 0.8000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.2500 0.0000 231.3500 0.8000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.2500 0.0000 227.3500 0.8000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.2500 0.0000 223.3500 0.8000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.2500 0.0000 219.3500 0.8000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.2500 0.0000 215.3500 0.8000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.2500 0.0000 211.3500 0.8000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.2500 0.0000 207.3500 0.8000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.2500 0.0000 203.3500 0.8000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.2500 0.0000 199.3500 0.8000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.2500 0.0000 195.3500 0.8000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.2500 0.0000 191.3500 0.8000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.2500 0.0000 187.3500 0.8000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.2500 0.0000 183.3500 0.8000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.2500 0.0000 179.3500 0.8000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.2500 0.0000 175.3500 0.8000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.2500 0.0000 171.3500 0.8000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.2500 0.0000 167.3500 0.8000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.2500 0.0000 163.3500 0.8000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.2500 0.0000 159.3500 0.8000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.2500 0.0000 155.3500 0.8000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.2500 0.0000 151.3500 0.8000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.2500 0.0000 147.3500 0.8000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.2500 0.0000 143.3500 0.8000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.2500 0.0000 139.3500 0.8000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.2500 0.0000 135.3500 0.8000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.2500 0.0000 131.3500 0.8000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.2500 0.0000 127.3500 0.8000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.2500 0.0000 123.3500 0.8000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.2500 0.0000 119.3500 0.8000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.2500 0.0000 115.3500 0.8000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.2500 0.0000 111.3500 0.8000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.2500 0.0000 107.3500 0.8000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.2500 0.0000 103.3500 0.8000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.2500 0.0000 99.3500 0.8000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.2500 0.0000 95.3500 0.8000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.2500 0.0000 91.3500 0.8000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.2500 0.0000 87.3500 0.8000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.2500 0.0000 83.3500 0.8000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.2500 0.0000 79.3500 0.8000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.2500 0.0000 75.3500 0.8000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.2500 0.0000 71.3500 0.8000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.2500 0.0000 67.3500 0.8000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.2500 0.0000 63.3500 0.8000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.2500 0.0000 59.3500 0.8000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.2500 0.0000 55.3500 0.8000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.2500 0.0000 51.3500 0.8000 ;
    END
  END D[0]
  PIN Q[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 687.2500 58.4000 687.3500 59.2000 ;
    END
  END Q[159]
  PIN Q[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 683.2500 58.4000 683.3500 59.2000 ;
    END
  END Q[158]
  PIN Q[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 679.2500 58.4000 679.3500 59.2000 ;
    END
  END Q[157]
  PIN Q[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 675.2500 58.4000 675.3500 59.2000 ;
    END
  END Q[156]
  PIN Q[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 671.2500 58.4000 671.3500 59.2000 ;
    END
  END Q[155]
  PIN Q[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 667.2500 58.4000 667.3500 59.2000 ;
    END
  END Q[154]
  PIN Q[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 663.2500 58.4000 663.3500 59.2000 ;
    END
  END Q[153]
  PIN Q[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 659.2500 58.4000 659.3500 59.2000 ;
    END
  END Q[152]
  PIN Q[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 655.2500 58.4000 655.3500 59.2000 ;
    END
  END Q[151]
  PIN Q[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 651.2500 58.4000 651.3500 59.2000 ;
    END
  END Q[150]
  PIN Q[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 647.2500 58.4000 647.3500 59.2000 ;
    END
  END Q[149]
  PIN Q[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 643.2500 58.4000 643.3500 59.2000 ;
    END
  END Q[148]
  PIN Q[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 639.2500 58.4000 639.3500 59.2000 ;
    END
  END Q[147]
  PIN Q[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 635.2500 58.4000 635.3500 59.2000 ;
    END
  END Q[146]
  PIN Q[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 631.2500 58.4000 631.3500 59.2000 ;
    END
  END Q[145]
  PIN Q[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 627.2500 58.4000 627.3500 59.2000 ;
    END
  END Q[144]
  PIN Q[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 623.2500 58.4000 623.3500 59.2000 ;
    END
  END Q[143]
  PIN Q[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 619.2500 58.4000 619.3500 59.2000 ;
    END
  END Q[142]
  PIN Q[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 615.2500 58.4000 615.3500 59.2000 ;
    END
  END Q[141]
  PIN Q[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 611.2500 58.4000 611.3500 59.2000 ;
    END
  END Q[140]
  PIN Q[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 607.2500 58.4000 607.3500 59.2000 ;
    END
  END Q[139]
  PIN Q[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 603.2500 58.4000 603.3500 59.2000 ;
    END
  END Q[138]
  PIN Q[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 599.2500 58.4000 599.3500 59.2000 ;
    END
  END Q[137]
  PIN Q[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 595.2500 58.4000 595.3500 59.2000 ;
    END
  END Q[136]
  PIN Q[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 591.2500 58.4000 591.3500 59.2000 ;
    END
  END Q[135]
  PIN Q[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 587.2500 58.4000 587.3500 59.2000 ;
    END
  END Q[134]
  PIN Q[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 583.2500 58.4000 583.3500 59.2000 ;
    END
  END Q[133]
  PIN Q[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 579.2500 58.4000 579.3500 59.2000 ;
    END
  END Q[132]
  PIN Q[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 575.2500 58.4000 575.3500 59.2000 ;
    END
  END Q[131]
  PIN Q[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 571.2500 58.4000 571.3500 59.2000 ;
    END
  END Q[130]
  PIN Q[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 567.2500 58.4000 567.3500 59.2000 ;
    END
  END Q[129]
  PIN Q[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 563.2500 58.4000 563.3500 59.2000 ;
    END
  END Q[128]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 559.2500 58.4000 559.3500 59.2000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 555.2500 58.4000 555.3500 59.2000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 551.2500 58.4000 551.3500 59.2000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 547.2500 58.4000 547.3500 59.2000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 543.2500 58.4000 543.3500 59.2000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 539.2500 58.4000 539.3500 59.2000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 535.2500 58.4000 535.3500 59.2000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 531.2500 58.4000 531.3500 59.2000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 527.2500 58.4000 527.3500 59.2000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 523.2500 58.4000 523.3500 59.2000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 519.2500 58.4000 519.3500 59.2000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 515.2500 58.4000 515.3500 59.2000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 511.2500 58.4000 511.3500 59.2000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 507.2500 58.4000 507.3500 59.2000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 503.2500 58.4000 503.3500 59.2000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 499.2500 58.4000 499.3500 59.2000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 495.2500 58.4000 495.3500 59.2000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 491.2500 58.4000 491.3500 59.2000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 487.2500 58.4000 487.3500 59.2000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 483.2500 58.4000 483.3500 59.2000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 479.2500 58.4000 479.3500 59.2000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 475.2500 58.4000 475.3500 59.2000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 471.2500 58.4000 471.3500 59.2000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 467.2500 58.4000 467.3500 59.2000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 463.2500 58.4000 463.3500 59.2000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 459.2500 58.4000 459.3500 59.2000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 455.2500 58.4000 455.3500 59.2000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 451.2500 58.4000 451.3500 59.2000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.2500 58.4000 447.3500 59.2000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.2500 58.4000 443.3500 59.2000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.2500 58.4000 439.3500 59.2000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.2500 58.4000 435.3500 59.2000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 431.2500 58.4000 431.3500 59.2000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.2500 58.4000 427.3500 59.2000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.2500 58.4000 423.3500 59.2000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.2500 58.4000 419.3500 59.2000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.2500 58.4000 415.3500 59.2000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 411.2500 58.4000 411.3500 59.2000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.2500 58.4000 407.3500 59.2000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.2500 58.4000 403.3500 59.2000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.2500 58.4000 399.3500 59.2000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.2500 58.4000 395.3500 59.2000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.2500 58.4000 391.3500 59.2000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.2500 58.4000 387.3500 59.2000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.2500 58.4000 383.3500 59.2000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 379.2500 58.4000 379.3500 59.2000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.2500 58.4000 375.3500 59.2000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.2500 58.4000 371.3500 59.2000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.2500 58.4000 367.3500 59.2000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.2500 58.4000 363.3500 59.2000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.2500 58.4000 359.3500 59.2000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.2500 58.4000 355.3500 59.2000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.2500 58.4000 351.3500 59.2000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.2500 58.4000 347.3500 59.2000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.2500 58.4000 343.3500 59.2000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.2500 58.4000 339.3500 59.2000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.2500 58.4000 335.3500 59.2000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.2500 58.4000 331.3500 59.2000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.2500 58.4000 327.3500 59.2000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.2500 58.4000 323.3500 59.2000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 319.2500 58.4000 319.3500 59.2000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.2500 58.4000 315.3500 59.2000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.2500 58.4000 311.3500 59.2000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 307.2500 58.4000 307.3500 59.2000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.2500 58.4000 303.3500 59.2000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 299.2500 58.4000 299.3500 59.2000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 295.2500 58.4000 295.3500 59.2000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.2500 58.4000 291.3500 59.2000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 287.2500 58.4000 287.3500 59.2000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 283.2500 58.4000 283.3500 59.2000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 279.2500 58.4000 279.3500 59.2000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 275.2500 58.4000 275.3500 59.2000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 271.2500 58.4000 271.3500 59.2000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.2500 58.4000 267.3500 59.2000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 263.2500 58.4000 263.3500 59.2000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.2500 58.4000 259.3500 59.2000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.2500 58.4000 255.3500 59.2000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 251.2500 58.4000 251.3500 59.2000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.2500 58.4000 247.3500 59.2000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.2500 58.4000 243.3500 59.2000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 239.2500 58.4000 239.3500 59.2000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.2500 58.4000 235.3500 59.2000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.2500 58.4000 231.3500 59.2000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.2500 58.4000 227.3500 59.2000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.2500 58.4000 223.3500 59.2000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.2500 58.4000 219.3500 59.2000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.2500 58.4000 215.3500 59.2000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.2500 58.4000 211.3500 59.2000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.2500 58.4000 207.3500 59.2000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.2500 58.4000 203.3500 59.2000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.2500 58.4000 199.3500 59.2000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.2500 58.4000 195.3500 59.2000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.2500 58.4000 191.3500 59.2000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.2500 58.4000 187.3500 59.2000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.2500 58.4000 183.3500 59.2000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.2500 58.4000 179.3500 59.2000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.2500 58.4000 175.3500 59.2000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.2500 58.4000 171.3500 59.2000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.2500 58.4000 167.3500 59.2000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.2500 58.4000 163.3500 59.2000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.2500 58.4000 159.3500 59.2000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.2500 58.4000 155.3500 59.2000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.2500 58.4000 151.3500 59.2000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.2500 58.4000 147.3500 59.2000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.2500 58.4000 143.3500 59.2000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.2500 58.4000 139.3500 59.2000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.2500 58.4000 135.3500 59.2000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.2500 58.4000 131.3500 59.2000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.2500 58.4000 127.3500 59.2000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.2500 58.4000 123.3500 59.2000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.2500 58.4000 119.3500 59.2000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.2500 58.4000 115.3500 59.2000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.2500 58.4000 111.3500 59.2000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.2500 58.4000 107.3500 59.2000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.2500 58.4000 103.3500 59.2000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.2500 58.4000 99.3500 59.2000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.2500 58.4000 95.3500 59.2000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.2500 58.4000 91.3500 59.2000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.2500 58.4000 87.3500 59.2000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.2500 58.4000 83.3500 59.2000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.2500 58.4000 79.3500 59.2000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.2500 58.4000 75.3500 59.2000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.2500 58.4000 71.3500 59.2000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.2500 58.4000 67.3500 59.2000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.2500 58.4000 63.3500 59.2000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.2500 58.4000 59.3500 59.2000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.2500 58.4000 55.3500 59.2000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.2500 58.4000 51.3500 59.2000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.3500 0.8000 19.4500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 39.3500 0.8000 39.4500 ;
    END
  END WEN
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 35.3500 0.8000 35.4500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 31.3500 0.8000 31.4500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.3500 0.8000 27.4500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 157.1100 8.0000 158.1100 51.2000 ;
        RECT 88.5550 8.0000 89.5550 51.2000 ;
        RECT 20.0000 8.0000 21.0000 51.2000 ;
        RECT 362.7750 8.0000 363.7750 51.2000 ;
        RECT 294.2200 8.0000 295.2200 51.2000 ;
        RECT 225.6650 8.0000 226.6650 51.2000 ;
        RECT 499.8850 8.0000 500.8850 51.2000 ;
        RECT 431.3300 8.0000 432.3300 51.2000 ;
        RECT 636.9950 8.0000 637.9950 51.2000 ;
        RECT 568.4400 8.0000 569.4400 51.2000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 159.1100 8.0000 160.1100 51.2000 ;
        RECT 90.5550 8.0000 91.5550 51.2000 ;
        RECT 22.0000 8.0000 23.0000 51.2000 ;
        RECT 364.7750 8.0000 365.7750 51.2000 ;
        RECT 296.2200 8.0000 297.2200 51.2000 ;
        RECT 227.6650 8.0000 228.6650 51.2000 ;
        RECT 501.8850 8.0000 502.8850 51.2000 ;
        RECT 433.3300 8.0000 434.3300 51.2000 ;
        RECT 638.9950 8.0000 639.9950 51.2000 ;
        RECT 570.4400 8.0000 571.4400 51.2000 ;
        RECT 22.0000 7.8350 23.0000 8.1650 ;
        RECT 90.5550 7.8350 91.5550 8.1650 ;
        RECT 159.1100 7.8350 160.1100 8.1650 ;
        RECT 227.6650 7.8350 228.6650 8.1650 ;
        RECT 296.2200 7.8350 297.2200 8.1650 ;
        RECT 364.7750 7.8350 365.7750 8.1650 ;
        RECT 433.3300 7.8350 434.3300 8.1650 ;
        RECT 501.8850 7.8350 502.8850 8.1650 ;
        RECT 570.4400 7.8350 571.4400 8.1650 ;
        RECT 638.9950 7.8350 639.9950 8.1650 ;
        RECT 22.0000 51.0350 23.0000 51.3650 ;
        RECT 90.5550 51.0350 91.5550 51.3650 ;
        RECT 159.1100 51.0350 160.1100 51.3650 ;
        RECT 227.6650 51.0350 228.6650 51.3650 ;
        RECT 296.2200 51.0350 297.2200 51.3650 ;
        RECT 364.7750 51.0350 365.7750 51.3650 ;
        RECT 433.3300 51.0350 434.3300 51.3650 ;
        RECT 501.8850 51.0350 502.8850 51.3650 ;
        RECT 570.4400 51.0350 571.4400 51.3650 ;
        RECT 638.9950 51.0350 639.9950 51.3650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 739.0000 59.2000 ;
    LAYER M2 ;
      RECT 687.4500 58.3000 739.0000 59.2000 ;
      RECT 683.4500 58.3000 687.1500 59.2000 ;
      RECT 679.4500 58.3000 683.1500 59.2000 ;
      RECT 675.4500 58.3000 679.1500 59.2000 ;
      RECT 671.4500 58.3000 675.1500 59.2000 ;
      RECT 667.4500 58.3000 671.1500 59.2000 ;
      RECT 663.4500 58.3000 667.1500 59.2000 ;
      RECT 659.4500 58.3000 663.1500 59.2000 ;
      RECT 655.4500 58.3000 659.1500 59.2000 ;
      RECT 651.4500 58.3000 655.1500 59.2000 ;
      RECT 647.4500 58.3000 651.1500 59.2000 ;
      RECT 643.4500 58.3000 647.1500 59.2000 ;
      RECT 639.4500 58.3000 643.1500 59.2000 ;
      RECT 635.4500 58.3000 639.1500 59.2000 ;
      RECT 631.4500 58.3000 635.1500 59.2000 ;
      RECT 627.4500 58.3000 631.1500 59.2000 ;
      RECT 623.4500 58.3000 627.1500 59.2000 ;
      RECT 619.4500 58.3000 623.1500 59.2000 ;
      RECT 615.4500 58.3000 619.1500 59.2000 ;
      RECT 611.4500 58.3000 615.1500 59.2000 ;
      RECT 607.4500 58.3000 611.1500 59.2000 ;
      RECT 603.4500 58.3000 607.1500 59.2000 ;
      RECT 599.4500 58.3000 603.1500 59.2000 ;
      RECT 595.4500 58.3000 599.1500 59.2000 ;
      RECT 591.4500 58.3000 595.1500 59.2000 ;
      RECT 587.4500 58.3000 591.1500 59.2000 ;
      RECT 583.4500 58.3000 587.1500 59.2000 ;
      RECT 579.4500 58.3000 583.1500 59.2000 ;
      RECT 575.4500 58.3000 579.1500 59.2000 ;
      RECT 571.4500 58.3000 575.1500 59.2000 ;
      RECT 567.4500 58.3000 571.1500 59.2000 ;
      RECT 563.4500 58.3000 567.1500 59.2000 ;
      RECT 559.4500 58.3000 563.1500 59.2000 ;
      RECT 555.4500 58.3000 559.1500 59.2000 ;
      RECT 551.4500 58.3000 555.1500 59.2000 ;
      RECT 547.4500 58.3000 551.1500 59.2000 ;
      RECT 543.4500 58.3000 547.1500 59.2000 ;
      RECT 539.4500 58.3000 543.1500 59.2000 ;
      RECT 535.4500 58.3000 539.1500 59.2000 ;
      RECT 531.4500 58.3000 535.1500 59.2000 ;
      RECT 527.4500 58.3000 531.1500 59.2000 ;
      RECT 523.4500 58.3000 527.1500 59.2000 ;
      RECT 519.4500 58.3000 523.1500 59.2000 ;
      RECT 515.4500 58.3000 519.1500 59.2000 ;
      RECT 511.4500 58.3000 515.1500 59.2000 ;
      RECT 507.4500 58.3000 511.1500 59.2000 ;
      RECT 503.4500 58.3000 507.1500 59.2000 ;
      RECT 499.4500 58.3000 503.1500 59.2000 ;
      RECT 495.4500 58.3000 499.1500 59.2000 ;
      RECT 491.4500 58.3000 495.1500 59.2000 ;
      RECT 487.4500 58.3000 491.1500 59.2000 ;
      RECT 483.4500 58.3000 487.1500 59.2000 ;
      RECT 479.4500 58.3000 483.1500 59.2000 ;
      RECT 475.4500 58.3000 479.1500 59.2000 ;
      RECT 471.4500 58.3000 475.1500 59.2000 ;
      RECT 467.4500 58.3000 471.1500 59.2000 ;
      RECT 463.4500 58.3000 467.1500 59.2000 ;
      RECT 459.4500 58.3000 463.1500 59.2000 ;
      RECT 455.4500 58.3000 459.1500 59.2000 ;
      RECT 451.4500 58.3000 455.1500 59.2000 ;
      RECT 447.4500 58.3000 451.1500 59.2000 ;
      RECT 443.4500 58.3000 447.1500 59.2000 ;
      RECT 439.4500 58.3000 443.1500 59.2000 ;
      RECT 435.4500 58.3000 439.1500 59.2000 ;
      RECT 431.4500 58.3000 435.1500 59.2000 ;
      RECT 427.4500 58.3000 431.1500 59.2000 ;
      RECT 423.4500 58.3000 427.1500 59.2000 ;
      RECT 419.4500 58.3000 423.1500 59.2000 ;
      RECT 415.4500 58.3000 419.1500 59.2000 ;
      RECT 411.4500 58.3000 415.1500 59.2000 ;
      RECT 407.4500 58.3000 411.1500 59.2000 ;
      RECT 403.4500 58.3000 407.1500 59.2000 ;
      RECT 399.4500 58.3000 403.1500 59.2000 ;
      RECT 395.4500 58.3000 399.1500 59.2000 ;
      RECT 391.4500 58.3000 395.1500 59.2000 ;
      RECT 387.4500 58.3000 391.1500 59.2000 ;
      RECT 383.4500 58.3000 387.1500 59.2000 ;
      RECT 379.4500 58.3000 383.1500 59.2000 ;
      RECT 375.4500 58.3000 379.1500 59.2000 ;
      RECT 371.4500 58.3000 375.1500 59.2000 ;
      RECT 367.4500 58.3000 371.1500 59.2000 ;
      RECT 363.4500 58.3000 367.1500 59.2000 ;
      RECT 359.4500 58.3000 363.1500 59.2000 ;
      RECT 355.4500 58.3000 359.1500 59.2000 ;
      RECT 351.4500 58.3000 355.1500 59.2000 ;
      RECT 347.4500 58.3000 351.1500 59.2000 ;
      RECT 343.4500 58.3000 347.1500 59.2000 ;
      RECT 339.4500 58.3000 343.1500 59.2000 ;
      RECT 335.4500 58.3000 339.1500 59.2000 ;
      RECT 331.4500 58.3000 335.1500 59.2000 ;
      RECT 327.4500 58.3000 331.1500 59.2000 ;
      RECT 323.4500 58.3000 327.1500 59.2000 ;
      RECT 319.4500 58.3000 323.1500 59.2000 ;
      RECT 315.4500 58.3000 319.1500 59.2000 ;
      RECT 311.4500 58.3000 315.1500 59.2000 ;
      RECT 307.4500 58.3000 311.1500 59.2000 ;
      RECT 303.4500 58.3000 307.1500 59.2000 ;
      RECT 299.4500 58.3000 303.1500 59.2000 ;
      RECT 295.4500 58.3000 299.1500 59.2000 ;
      RECT 291.4500 58.3000 295.1500 59.2000 ;
      RECT 287.4500 58.3000 291.1500 59.2000 ;
      RECT 283.4500 58.3000 287.1500 59.2000 ;
      RECT 279.4500 58.3000 283.1500 59.2000 ;
      RECT 275.4500 58.3000 279.1500 59.2000 ;
      RECT 271.4500 58.3000 275.1500 59.2000 ;
      RECT 267.4500 58.3000 271.1500 59.2000 ;
      RECT 263.4500 58.3000 267.1500 59.2000 ;
      RECT 259.4500 58.3000 263.1500 59.2000 ;
      RECT 255.4500 58.3000 259.1500 59.2000 ;
      RECT 251.4500 58.3000 255.1500 59.2000 ;
      RECT 247.4500 58.3000 251.1500 59.2000 ;
      RECT 243.4500 58.3000 247.1500 59.2000 ;
      RECT 239.4500 58.3000 243.1500 59.2000 ;
      RECT 235.4500 58.3000 239.1500 59.2000 ;
      RECT 231.4500 58.3000 235.1500 59.2000 ;
      RECT 227.4500 58.3000 231.1500 59.2000 ;
      RECT 223.4500 58.3000 227.1500 59.2000 ;
      RECT 219.4500 58.3000 223.1500 59.2000 ;
      RECT 215.4500 58.3000 219.1500 59.2000 ;
      RECT 211.4500 58.3000 215.1500 59.2000 ;
      RECT 207.4500 58.3000 211.1500 59.2000 ;
      RECT 203.4500 58.3000 207.1500 59.2000 ;
      RECT 199.4500 58.3000 203.1500 59.2000 ;
      RECT 195.4500 58.3000 199.1500 59.2000 ;
      RECT 191.4500 58.3000 195.1500 59.2000 ;
      RECT 187.4500 58.3000 191.1500 59.2000 ;
      RECT 183.4500 58.3000 187.1500 59.2000 ;
      RECT 179.4500 58.3000 183.1500 59.2000 ;
      RECT 175.4500 58.3000 179.1500 59.2000 ;
      RECT 171.4500 58.3000 175.1500 59.2000 ;
      RECT 167.4500 58.3000 171.1500 59.2000 ;
      RECT 163.4500 58.3000 167.1500 59.2000 ;
      RECT 159.4500 58.3000 163.1500 59.2000 ;
      RECT 155.4500 58.3000 159.1500 59.2000 ;
      RECT 151.4500 58.3000 155.1500 59.2000 ;
      RECT 147.4500 58.3000 151.1500 59.2000 ;
      RECT 143.4500 58.3000 147.1500 59.2000 ;
      RECT 139.4500 58.3000 143.1500 59.2000 ;
      RECT 135.4500 58.3000 139.1500 59.2000 ;
      RECT 131.4500 58.3000 135.1500 59.2000 ;
      RECT 127.4500 58.3000 131.1500 59.2000 ;
      RECT 123.4500 58.3000 127.1500 59.2000 ;
      RECT 119.4500 58.3000 123.1500 59.2000 ;
      RECT 115.4500 58.3000 119.1500 59.2000 ;
      RECT 111.4500 58.3000 115.1500 59.2000 ;
      RECT 107.4500 58.3000 111.1500 59.2000 ;
      RECT 103.4500 58.3000 107.1500 59.2000 ;
      RECT 99.4500 58.3000 103.1500 59.2000 ;
      RECT 95.4500 58.3000 99.1500 59.2000 ;
      RECT 91.4500 58.3000 95.1500 59.2000 ;
      RECT 87.4500 58.3000 91.1500 59.2000 ;
      RECT 83.4500 58.3000 87.1500 59.2000 ;
      RECT 79.4500 58.3000 83.1500 59.2000 ;
      RECT 75.4500 58.3000 79.1500 59.2000 ;
      RECT 71.4500 58.3000 75.1500 59.2000 ;
      RECT 67.4500 58.3000 71.1500 59.2000 ;
      RECT 63.4500 58.3000 67.1500 59.2000 ;
      RECT 59.4500 58.3000 63.1500 59.2000 ;
      RECT 55.4500 58.3000 59.1500 59.2000 ;
      RECT 51.4500 58.3000 55.1500 59.2000 ;
      RECT 0.0000 58.3000 51.1500 59.2000 ;
      RECT 0.0000 0.9000 739.0000 58.3000 ;
      RECT 687.4500 0.0000 739.0000 0.9000 ;
      RECT 683.4500 0.0000 687.1500 0.9000 ;
      RECT 679.4500 0.0000 683.1500 0.9000 ;
      RECT 675.4500 0.0000 679.1500 0.9000 ;
      RECT 671.4500 0.0000 675.1500 0.9000 ;
      RECT 667.4500 0.0000 671.1500 0.9000 ;
      RECT 663.4500 0.0000 667.1500 0.9000 ;
      RECT 659.4500 0.0000 663.1500 0.9000 ;
      RECT 655.4500 0.0000 659.1500 0.9000 ;
      RECT 651.4500 0.0000 655.1500 0.9000 ;
      RECT 647.4500 0.0000 651.1500 0.9000 ;
      RECT 643.4500 0.0000 647.1500 0.9000 ;
      RECT 639.4500 0.0000 643.1500 0.9000 ;
      RECT 635.4500 0.0000 639.1500 0.9000 ;
      RECT 631.4500 0.0000 635.1500 0.9000 ;
      RECT 627.4500 0.0000 631.1500 0.9000 ;
      RECT 623.4500 0.0000 627.1500 0.9000 ;
      RECT 619.4500 0.0000 623.1500 0.9000 ;
      RECT 615.4500 0.0000 619.1500 0.9000 ;
      RECT 611.4500 0.0000 615.1500 0.9000 ;
      RECT 607.4500 0.0000 611.1500 0.9000 ;
      RECT 603.4500 0.0000 607.1500 0.9000 ;
      RECT 599.4500 0.0000 603.1500 0.9000 ;
      RECT 595.4500 0.0000 599.1500 0.9000 ;
      RECT 591.4500 0.0000 595.1500 0.9000 ;
      RECT 587.4500 0.0000 591.1500 0.9000 ;
      RECT 583.4500 0.0000 587.1500 0.9000 ;
      RECT 579.4500 0.0000 583.1500 0.9000 ;
      RECT 575.4500 0.0000 579.1500 0.9000 ;
      RECT 571.4500 0.0000 575.1500 0.9000 ;
      RECT 567.4500 0.0000 571.1500 0.9000 ;
      RECT 563.4500 0.0000 567.1500 0.9000 ;
      RECT 559.4500 0.0000 563.1500 0.9000 ;
      RECT 555.4500 0.0000 559.1500 0.9000 ;
      RECT 551.4500 0.0000 555.1500 0.9000 ;
      RECT 547.4500 0.0000 551.1500 0.9000 ;
      RECT 543.4500 0.0000 547.1500 0.9000 ;
      RECT 539.4500 0.0000 543.1500 0.9000 ;
      RECT 535.4500 0.0000 539.1500 0.9000 ;
      RECT 531.4500 0.0000 535.1500 0.9000 ;
      RECT 527.4500 0.0000 531.1500 0.9000 ;
      RECT 523.4500 0.0000 527.1500 0.9000 ;
      RECT 519.4500 0.0000 523.1500 0.9000 ;
      RECT 515.4500 0.0000 519.1500 0.9000 ;
      RECT 511.4500 0.0000 515.1500 0.9000 ;
      RECT 507.4500 0.0000 511.1500 0.9000 ;
      RECT 503.4500 0.0000 507.1500 0.9000 ;
      RECT 499.4500 0.0000 503.1500 0.9000 ;
      RECT 495.4500 0.0000 499.1500 0.9000 ;
      RECT 491.4500 0.0000 495.1500 0.9000 ;
      RECT 487.4500 0.0000 491.1500 0.9000 ;
      RECT 483.4500 0.0000 487.1500 0.9000 ;
      RECT 479.4500 0.0000 483.1500 0.9000 ;
      RECT 475.4500 0.0000 479.1500 0.9000 ;
      RECT 471.4500 0.0000 475.1500 0.9000 ;
      RECT 467.4500 0.0000 471.1500 0.9000 ;
      RECT 463.4500 0.0000 467.1500 0.9000 ;
      RECT 459.4500 0.0000 463.1500 0.9000 ;
      RECT 455.4500 0.0000 459.1500 0.9000 ;
      RECT 451.4500 0.0000 455.1500 0.9000 ;
      RECT 447.4500 0.0000 451.1500 0.9000 ;
      RECT 443.4500 0.0000 447.1500 0.9000 ;
      RECT 439.4500 0.0000 443.1500 0.9000 ;
      RECT 435.4500 0.0000 439.1500 0.9000 ;
      RECT 431.4500 0.0000 435.1500 0.9000 ;
      RECT 427.4500 0.0000 431.1500 0.9000 ;
      RECT 423.4500 0.0000 427.1500 0.9000 ;
      RECT 419.4500 0.0000 423.1500 0.9000 ;
      RECT 415.4500 0.0000 419.1500 0.9000 ;
      RECT 411.4500 0.0000 415.1500 0.9000 ;
      RECT 407.4500 0.0000 411.1500 0.9000 ;
      RECT 403.4500 0.0000 407.1500 0.9000 ;
      RECT 399.4500 0.0000 403.1500 0.9000 ;
      RECT 395.4500 0.0000 399.1500 0.9000 ;
      RECT 391.4500 0.0000 395.1500 0.9000 ;
      RECT 387.4500 0.0000 391.1500 0.9000 ;
      RECT 383.4500 0.0000 387.1500 0.9000 ;
      RECT 379.4500 0.0000 383.1500 0.9000 ;
      RECT 375.4500 0.0000 379.1500 0.9000 ;
      RECT 371.4500 0.0000 375.1500 0.9000 ;
      RECT 367.4500 0.0000 371.1500 0.9000 ;
      RECT 363.4500 0.0000 367.1500 0.9000 ;
      RECT 359.4500 0.0000 363.1500 0.9000 ;
      RECT 355.4500 0.0000 359.1500 0.9000 ;
      RECT 351.4500 0.0000 355.1500 0.9000 ;
      RECT 347.4500 0.0000 351.1500 0.9000 ;
      RECT 343.4500 0.0000 347.1500 0.9000 ;
      RECT 339.4500 0.0000 343.1500 0.9000 ;
      RECT 335.4500 0.0000 339.1500 0.9000 ;
      RECT 331.4500 0.0000 335.1500 0.9000 ;
      RECT 327.4500 0.0000 331.1500 0.9000 ;
      RECT 323.4500 0.0000 327.1500 0.9000 ;
      RECT 319.4500 0.0000 323.1500 0.9000 ;
      RECT 315.4500 0.0000 319.1500 0.9000 ;
      RECT 311.4500 0.0000 315.1500 0.9000 ;
      RECT 307.4500 0.0000 311.1500 0.9000 ;
      RECT 303.4500 0.0000 307.1500 0.9000 ;
      RECT 299.4500 0.0000 303.1500 0.9000 ;
      RECT 295.4500 0.0000 299.1500 0.9000 ;
      RECT 291.4500 0.0000 295.1500 0.9000 ;
      RECT 287.4500 0.0000 291.1500 0.9000 ;
      RECT 283.4500 0.0000 287.1500 0.9000 ;
      RECT 279.4500 0.0000 283.1500 0.9000 ;
      RECT 275.4500 0.0000 279.1500 0.9000 ;
      RECT 271.4500 0.0000 275.1500 0.9000 ;
      RECT 267.4500 0.0000 271.1500 0.9000 ;
      RECT 263.4500 0.0000 267.1500 0.9000 ;
      RECT 259.4500 0.0000 263.1500 0.9000 ;
      RECT 255.4500 0.0000 259.1500 0.9000 ;
      RECT 251.4500 0.0000 255.1500 0.9000 ;
      RECT 247.4500 0.0000 251.1500 0.9000 ;
      RECT 243.4500 0.0000 247.1500 0.9000 ;
      RECT 239.4500 0.0000 243.1500 0.9000 ;
      RECT 235.4500 0.0000 239.1500 0.9000 ;
      RECT 231.4500 0.0000 235.1500 0.9000 ;
      RECT 227.4500 0.0000 231.1500 0.9000 ;
      RECT 223.4500 0.0000 227.1500 0.9000 ;
      RECT 219.4500 0.0000 223.1500 0.9000 ;
      RECT 215.4500 0.0000 219.1500 0.9000 ;
      RECT 211.4500 0.0000 215.1500 0.9000 ;
      RECT 207.4500 0.0000 211.1500 0.9000 ;
      RECT 203.4500 0.0000 207.1500 0.9000 ;
      RECT 199.4500 0.0000 203.1500 0.9000 ;
      RECT 195.4500 0.0000 199.1500 0.9000 ;
      RECT 191.4500 0.0000 195.1500 0.9000 ;
      RECT 187.4500 0.0000 191.1500 0.9000 ;
      RECT 183.4500 0.0000 187.1500 0.9000 ;
      RECT 179.4500 0.0000 183.1500 0.9000 ;
      RECT 175.4500 0.0000 179.1500 0.9000 ;
      RECT 171.4500 0.0000 175.1500 0.9000 ;
      RECT 167.4500 0.0000 171.1500 0.9000 ;
      RECT 163.4500 0.0000 167.1500 0.9000 ;
      RECT 159.4500 0.0000 163.1500 0.9000 ;
      RECT 155.4500 0.0000 159.1500 0.9000 ;
      RECT 151.4500 0.0000 155.1500 0.9000 ;
      RECT 147.4500 0.0000 151.1500 0.9000 ;
      RECT 143.4500 0.0000 147.1500 0.9000 ;
      RECT 139.4500 0.0000 143.1500 0.9000 ;
      RECT 135.4500 0.0000 139.1500 0.9000 ;
      RECT 131.4500 0.0000 135.1500 0.9000 ;
      RECT 127.4500 0.0000 131.1500 0.9000 ;
      RECT 123.4500 0.0000 127.1500 0.9000 ;
      RECT 119.4500 0.0000 123.1500 0.9000 ;
      RECT 115.4500 0.0000 119.1500 0.9000 ;
      RECT 111.4500 0.0000 115.1500 0.9000 ;
      RECT 107.4500 0.0000 111.1500 0.9000 ;
      RECT 103.4500 0.0000 107.1500 0.9000 ;
      RECT 99.4500 0.0000 103.1500 0.9000 ;
      RECT 95.4500 0.0000 99.1500 0.9000 ;
      RECT 91.4500 0.0000 95.1500 0.9000 ;
      RECT 87.4500 0.0000 91.1500 0.9000 ;
      RECT 83.4500 0.0000 87.1500 0.9000 ;
      RECT 79.4500 0.0000 83.1500 0.9000 ;
      RECT 75.4500 0.0000 79.1500 0.9000 ;
      RECT 71.4500 0.0000 75.1500 0.9000 ;
      RECT 67.4500 0.0000 71.1500 0.9000 ;
      RECT 63.4500 0.0000 67.1500 0.9000 ;
      RECT 59.4500 0.0000 63.1500 0.9000 ;
      RECT 55.4500 0.0000 59.1500 0.9000 ;
      RECT 51.4500 0.0000 55.1500 0.9000 ;
      RECT 0.0000 0.0000 51.1500 0.9000 ;
    LAYER M3 ;
      RECT 0.0000 39.5500 739.0000 59.2000 ;
      RECT 0.9000 39.2500 739.0000 39.5500 ;
      RECT 0.0000 35.5500 739.0000 39.2500 ;
      RECT 0.9000 35.2500 739.0000 35.5500 ;
      RECT 0.0000 31.5500 739.0000 35.2500 ;
      RECT 0.9000 31.2500 739.0000 31.5500 ;
      RECT 0.0000 27.5500 739.0000 31.2500 ;
      RECT 0.9000 27.2500 739.0000 27.5500 ;
      RECT 0.0000 23.5500 739.0000 27.2500 ;
      RECT 0.9000 23.2500 739.0000 23.5500 ;
      RECT 0.0000 19.5500 739.0000 23.2500 ;
      RECT 0.9000 19.2500 739.0000 19.5500 ;
      RECT 0.0000 0.0000 739.0000 19.2500 ;
    LAYER M4 ;
      RECT 0.0000 51.5250 739.0000 59.2000 ;
      RECT 571.6000 51.3600 638.8350 51.5250 ;
      RECT 503.0450 51.3600 570.2800 51.5250 ;
      RECT 434.4900 51.3600 501.7250 51.5250 ;
      RECT 365.9350 51.3600 433.1700 51.5250 ;
      RECT 297.3800 51.3600 364.6150 51.5250 ;
      RECT 228.8250 51.3600 296.0600 51.5250 ;
      RECT 160.2700 51.3600 227.5050 51.5250 ;
      RECT 91.7150 51.3600 158.9500 51.5250 ;
      RECT 23.1600 51.3600 90.3950 51.5250 ;
      RECT 0.0000 51.3600 21.8400 51.5250 ;
      RECT 638.1550 7.8400 638.8350 51.3600 ;
      RECT 571.6000 7.8400 636.8350 51.3600 ;
      RECT 569.6000 7.8400 570.2800 51.3600 ;
      RECT 503.0450 7.8400 568.2800 51.3600 ;
      RECT 501.0450 7.8400 501.7250 51.3600 ;
      RECT 434.4900 7.8400 499.7250 51.3600 ;
      RECT 432.4900 7.8400 433.1700 51.3600 ;
      RECT 365.9350 7.8400 431.1700 51.3600 ;
      RECT 363.9350 7.8400 364.6150 51.3600 ;
      RECT 297.3800 7.8400 362.6150 51.3600 ;
      RECT 295.3800 7.8400 296.0600 51.3600 ;
      RECT 228.8250 7.8400 294.0600 51.3600 ;
      RECT 226.8250 7.8400 227.5050 51.3600 ;
      RECT 160.2700 7.8400 225.5050 51.3600 ;
      RECT 158.2700 7.8400 158.9500 51.3600 ;
      RECT 91.7150 7.8400 156.9500 51.3600 ;
      RECT 89.7150 7.8400 90.3950 51.3600 ;
      RECT 23.1600 7.8400 88.3950 51.3600 ;
      RECT 21.1600 7.8400 21.8400 51.3600 ;
      RECT 0.0000 7.8400 19.8400 51.3600 ;
      RECT 640.1550 7.6750 739.0000 51.5250 ;
      RECT 571.6000 7.6750 638.8350 7.8400 ;
      RECT 503.0450 7.6750 570.2800 7.8400 ;
      RECT 434.4900 7.6750 501.7250 7.8400 ;
      RECT 365.9350 7.6750 433.1700 7.8400 ;
      RECT 297.3800 7.6750 364.6150 7.8400 ;
      RECT 228.8250 7.6750 296.0600 7.8400 ;
      RECT 160.2700 7.6750 227.5050 7.8400 ;
      RECT 91.7150 7.6750 158.9500 7.8400 ;
      RECT 23.1600 7.6750 90.3950 7.8400 ;
      RECT 0.0000 7.6750 21.8400 7.8400 ;
      RECT 0.0000 0.0000 739.0000 7.6750 ;
  END
END sram_w16_2

END LIBRARY
